
module mux21_generic_n4_7 ( a, b, sel, y );
  input [3:0] a;
  input [3:0] b;
  output [3:0] y;
  input sel;


  mux21_28 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(sel), .y(y[0]) );
  mux21_27 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(sel), .y(y[1]) );
  mux21_26 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(sel), .y(y[2]) );
  mux21_25 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(sel), .y(y[3]) );
endmodule


module mux21_generic_n4_6 ( a, b, sel, y );
  input [3:0] a;
  input [3:0] b;
  output [3:0] y;
  input sel;


  mux21_24 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(sel), .y(y[0]) );
  mux21_23 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(sel), .y(y[1]) );
  mux21_22 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(sel), .y(y[2]) );
  mux21_21 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(sel), .y(y[3]) );
endmodule


module mux21_generic_n4_5 ( a, b, sel, y );
  input [3:0] a;
  input [3:0] b;
  output [3:0] y;
  input sel;


  mux21_20 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(sel), .y(y[0]) );
  mux21_19 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(sel), .y(y[1]) );
  mux21_18 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(sel), .y(y[2]) );
  mux21_17 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(sel), .y(y[3]) );
endmodule


module mux21_generic_n4_4 ( a, b, sel, y );
  input [3:0] a;
  input [3:0] b;
  output [3:0] y;
  input sel;


  mux21_16 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(sel), .y(y[0]) );
  mux21_15 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(sel), .y(y[1]) );
  mux21_14 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(sel), .y(y[2]) );
  mux21_13 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(sel), .y(y[3]) );
endmodule


module mux21_generic_n4_3 ( a, b, sel, y );
  input [3:0] a;
  input [3:0] b;
  output [3:0] y;
  input sel;


  mux21_12 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(sel), .y(y[0]) );
  mux21_11 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(sel), .y(y[1]) );
  mux21_10 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(sel), .y(y[2]) );
  mux21_9 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(sel), .y(y[3]) );
endmodule


module mux21_generic_n4_2 ( a, b, sel, y );
  input [3:0] a;
  input [3:0] b;
  output [3:0] y;
  input sel;


  mux21_8 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(sel), .y(y[0]) );
  mux21_7 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(sel), .y(y[1]) );
  mux21_6 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(sel), .y(y[2]) );
  mux21_5 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(sel), .y(y[3]) );
endmodule


module mux21_generic_n4_1 ( a, b, sel, y );
  input [3:0] a;
  input [3:0] b;
  output [3:0] y;
  input sel;


  mux21_4 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(sel), .y(y[0]) );
  mux21_3 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(sel), .y(y[1]) );
  mux21_2 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(sel), .y(y[2]) );
  mux21_1 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(sel), .y(y[3]) );
endmodule


module rca_n_n4_15 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_60 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_59 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_58 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_57 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_14 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_56 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_55 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_54 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_53 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_13 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_52 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_51 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_50 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_49 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_12 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_48 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_47 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_46 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_45 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_11 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_44 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_43 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_42 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_41 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_10 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_40 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_39 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_38 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_37 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_9 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_36 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_35 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_34 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_33 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_8 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_32 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_31 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_30 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_29 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_7 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_28 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_27 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_26 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_25 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_6 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_24 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_23 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_22 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_21 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_5 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_20 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_19 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_18 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_17 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_4 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_16 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_15 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_14 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_13 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_3 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_12 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_11 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_10 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_9 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_2 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_8 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_7 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_6 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_5 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module rca_n_n4_1 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_4 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_3 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_2 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_1 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module PG_31 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_223 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_159 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_30 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_222 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_158 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_29 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_221 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_157 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_28 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_220 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_156 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_27 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_219 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_155 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_26 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_218 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_154 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_25 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_217 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_153 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_24 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_216 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_152 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_23 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_215 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_151 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_22 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_214 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_150 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_21 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_213 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_149 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_20 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_212 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_148 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_19 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_211 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_147 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_18 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_210 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_146 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_17 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_209 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_145 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_16 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_208 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_144 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_15 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_207 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_143 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_14 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_206 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_142 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_13 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_205 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_141 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_12 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_204 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_140 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_11 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_203 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_139 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_10 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_202 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_138 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_9 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_201 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_137 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_8 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_200 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_136 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_7 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_199 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_135 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_6 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_198 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_134 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_5 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_197 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_133 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_4 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_196 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_132 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_3 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_195 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_131 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_2 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_194 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_130 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module PG_1 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_193 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_129 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module carry_select_block_n4_7 ( a, b, cin, s );
  input [3:0] a;
  input [3:0] b;
  output [3:0] s;
  input cin;

  wire   [3:0] sum_first_rca;
  wire   [3:0] sum_second_rca;

  rca_n_n4_14 first_rca ( .a(a), .b(b), .c_in(1'b0), .sum(sum_first_rca) );
  rca_n_n4_13 second_rca ( .a(a), .b(b), .c_in(1'b1), .sum(sum_second_rca) );
  mux21_generic_n4_7 mux ( .a(sum_first_rca), .b(sum_second_rca), .sel(cin), 
        .y(s) );
endmodule


module carry_select_block_n4_6 ( a, b, cin, s );
  input [3:0] a;
  input [3:0] b;
  output [3:0] s;
  input cin;

  wire   [3:0] sum_first_rca;
  wire   [3:0] sum_second_rca;

  rca_n_n4_12 first_rca ( .a(a), .b(b), .c_in(1'b0), .sum(sum_first_rca) );
  rca_n_n4_11 second_rca ( .a(a), .b(b), .c_in(1'b1), .sum(sum_second_rca) );
  mux21_generic_n4_6 mux ( .a(sum_first_rca), .b(sum_second_rca), .sel(cin), 
        .y(s) );
endmodule


module carry_select_block_n4_5 ( a, b, cin, s );
  input [3:0] a;
  input [3:0] b;
  output [3:0] s;
  input cin;

  wire   [3:0] sum_first_rca;
  wire   [3:0] sum_second_rca;

  rca_n_n4_10 first_rca ( .a(a), .b(b), .c_in(1'b0), .sum(sum_first_rca) );
  rca_n_n4_9 second_rca ( .a(a), .b(b), .c_in(1'b1), .sum(sum_second_rca) );
  mux21_generic_n4_5 mux ( .a(sum_first_rca), .b(sum_second_rca), .sel(cin), 
        .y(s) );
endmodule


module carry_select_block_n4_4 ( a, b, cin, s );
  input [3:0] a;
  input [3:0] b;
  output [3:0] s;
  input cin;

  wire   [3:0] sum_first_rca;
  wire   [3:0] sum_second_rca;

  rca_n_n4_8 first_rca ( .a(a), .b(b), .c_in(1'b0), .sum(sum_first_rca) );
  rca_n_n4_7 second_rca ( .a(a), .b(b), .c_in(1'b1), .sum(sum_second_rca) );
  mux21_generic_n4_4 mux ( .a(sum_first_rca), .b(sum_second_rca), .sel(cin), 
        .y(s) );
endmodule


module carry_select_block_n4_3 ( a, b, cin, s );
  input [3:0] a;
  input [3:0] b;
  output [3:0] s;
  input cin;

  wire   [3:0] sum_first_rca;
  wire   [3:0] sum_second_rca;

  rca_n_n4_6 first_rca ( .a(a), .b(b), .c_in(1'b0), .sum(sum_first_rca) );
  rca_n_n4_5 second_rca ( .a(a), .b(b), .c_in(1'b1), .sum(sum_second_rca) );
  mux21_generic_n4_3 mux ( .a(sum_first_rca), .b(sum_second_rca), .sel(cin), 
        .y(s) );
endmodule


module carry_select_block_n4_2 ( a, b, cin, s );
  input [3:0] a;
  input [3:0] b;
  output [3:0] s;
  input cin;

  wire   [3:0] sum_first_rca;
  wire   [3:0] sum_second_rca;

  rca_n_n4_4 first_rca ( .a(a), .b(b), .c_in(1'b0), .sum(sum_first_rca) );
  rca_n_n4_3 second_rca ( .a(a), .b(b), .c_in(1'b1), .sum(sum_second_rca) );
  mux21_generic_n4_2 mux ( .a(sum_first_rca), .b(sum_second_rca), .sel(cin), 
        .y(s) );
endmodule


module carry_select_block_n4_1 ( a, b, cin, s );
  input [3:0] a;
  input [3:0] b;
  output [3:0] s;
  input cin;

  wire   [3:0] sum_first_rca;
  wire   [3:0] sum_second_rca;

  rca_n_n4_2 first_rca ( .a(a), .b(b), .c_in(1'b0), .sum(sum_first_rca) );
  rca_n_n4_1 second_rca ( .a(a), .b(b), .c_in(1'b1), .sum(sum_second_rca) );
  mux21_generic_n4_1 mux ( .a(sum_first_rca), .b(sum_second_rca), .sel(cin), 
        .y(s) );
endmodule


module PG_general_26 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_412 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_194 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_411 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_25 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_410 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_193 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_409 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_24 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_408 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_192 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_407 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_23 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_406 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_191 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_405 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_22 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_404 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_190 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_403 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_21 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_402 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_189 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_401 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_20 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_400 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_188 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_399 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_19 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_398 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_187 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_397 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_18 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_396 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_186 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_395 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_17 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_394 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_185 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_393 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_16 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_392 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_184 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_391 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_15 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_390 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_183 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_389 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_14 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_388 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_182 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_387 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_13 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_386 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_181 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_385 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_12 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_383 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_179 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_382 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_11 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_381 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_178 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_380 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_10 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_379 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_177 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_378 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_9 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_377 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_176 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_376 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_8 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_375 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_175 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_374 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_7 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_373 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_174 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_372 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_6 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_371 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_173 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_370 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_5 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_368 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_171 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_367 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_4 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_366 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_170 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_365 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_3 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_364 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_169 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_363 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_2 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_360 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_166 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_359 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module PG_general_1 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_358 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_165 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_357 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module G_general_8 ( gkminj, gik, pik, gij );
  input gkminj, gik, pik;
  output gij;
  wire   and_out;

  and_2_384 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_180 or_gen ( .a(gik), .b(and_out), .y(gij) );
endmodule


module G_general_7 ( gkminj, gik, pik, gij );
  input gkminj, gik, pik;
  output gij;
  wire   and_out;

  and_2_369 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_172 or_gen ( .a(gik), .b(and_out), .y(gij) );
endmodule


module G_general_6 ( gkminj, gik, pik, gij );
  input gkminj, gik, pik;
  output gij;
  wire   and_out;

  and_2_362 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_168 or_gen ( .a(gik), .b(and_out), .y(gij) );
endmodule


module G_general_5 ( gkminj, gik, pik, gij );
  input gkminj, gik, pik;
  output gij;
  wire   and_out;

  and_2_361 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_167 or_gen ( .a(gik), .b(and_out), .y(gij) );
endmodule


module G_general_4 ( gkminj, gik, pik, gij );
  input gkminj, gik, pik;
  output gij;
  wire   and_out;

  and_2_356 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_164 or_gen ( .a(gik), .b(and_out), .y(gij) );
endmodule


module G_general_3 ( gkminj, gik, pik, gij );
  input gkminj, gik, pik;
  output gij;
  wire   and_out;

  and_2_355 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_163 or_gen ( .a(gik), .b(and_out), .y(gij) );
endmodule


module G_general_2 ( gkminj, gik, pik, gij );
  input gkminj, gik, pik;
  output gij;
  wire   and_out;

  and_2_354 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_162 or_gen ( .a(gik), .b(and_out), .y(gij) );
endmodule


module G_general_1 ( gkminj, gik, pik, gij );
  input gkminj, gik, pik;
  output gij;
  wire   and_out;

  and_2_353 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_161 or_gen ( .a(gik), .b(and_out), .y(gij) );
endmodule


module logic_31 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n4, n7, n8, n9;

  OAI22_X1 U1 ( .A1(n9), .A2(n4), .B1(r2), .B2(n8), .ZN(y) );
  AOI22_X1 U2 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U4 ( .A(r1), .ZN(n7) );
  INV_X1 U5 ( .A(r2), .ZN(n4) );
endmodule


module logic_30 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n4, n7, n8, n9;

  OAI22_X1 U1 ( .A1(n9), .A2(n4), .B1(r2), .B2(n8), .ZN(y) );
  AOI22_X1 U2 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U4 ( .A(r1), .ZN(n7) );
  INV_X1 U5 ( .A(r2), .ZN(n4) );
endmodule


module logic_29 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n4, n7, n8, n9;

  OAI22_X1 U1 ( .A1(n9), .A2(n4), .B1(r2), .B2(n8), .ZN(y) );
  AOI22_X1 U2 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U4 ( .A(r1), .ZN(n7) );
  INV_X1 U5 ( .A(r2), .ZN(n4) );
endmodule


module logic_28 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n4, n7, n8, n9;

  OAI22_X1 U1 ( .A1(n9), .A2(n4), .B1(r2), .B2(n8), .ZN(y) );
  AOI22_X1 U2 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U4 ( .A(r1), .ZN(n7) );
  INV_X1 U5 ( .A(r2), .ZN(n4) );
endmodule


module logic_27 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_26 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_25 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_24 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_23 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_22 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_21 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_20 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_19 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_18 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_17 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_16 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_15 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_14 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_13 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_12 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_11 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_10 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_9 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_8 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_7 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_6 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_5 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_4 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_3 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_2 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module logic_1 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n7, n8, n9, n10;

  OAI22_X1 U1 ( .A1(n10), .A2(n9), .B1(r2), .B2(n8), .ZN(y) );
  INV_X1 U2 ( .A(r2), .ZN(n9) );
  AOI22_X1 U3 ( .A1(s1), .A2(n7), .B1(s3), .B2(r1), .ZN(n10) );
  AOI22_X1 U4 ( .A1(s0), .A2(n7), .B1(s2), .B2(r1), .ZN(n8) );
  INV_X1 U5 ( .A(r1), .ZN(n7) );
endmodule


module not_n_n32_1 ( a, y );
  input [31:0] a;
  output [31:0] y;


  not_1_64 not_1_component_0 ( .a(a[0]), .y(y[0]) );
  not_1_63 not_1_component_1 ( .a(a[1]), .y(y[1]) );
  not_1_62 not_1_component_2 ( .a(a[2]), .y(y[2]) );
  not_1_61 not_1_component_3 ( .a(a[3]), .y(y[3]) );
  not_1_60 not_1_component_4 ( .a(a[4]), .y(y[4]) );
  not_1_59 not_1_component_5 ( .a(a[5]), .y(y[5]) );
  not_1_58 not_1_component_6 ( .a(a[6]), .y(y[6]) );
  not_1_57 not_1_component_7 ( .a(a[7]), .y(y[7]) );
  not_1_56 not_1_component_8 ( .a(a[8]), .y(y[8]) );
  not_1_55 not_1_component_9 ( .a(a[9]), .y(y[9]) );
  not_1_54 not_1_component_10 ( .a(a[10]), .y(y[10]) );
  not_1_53 not_1_component_11 ( .a(a[11]), .y(y[11]) );
  not_1_52 not_1_component_12 ( .a(a[12]), .y(y[12]) );
  not_1_51 not_1_component_13 ( .a(a[13]), .y(y[13]) );
  not_1_50 not_1_component_14 ( .a(a[14]), .y(y[14]) );
  not_1_49 not_1_component_15 ( .a(a[15]), .y(y[15]) );
  not_1_48 not_1_component_16 ( .a(a[16]), .y(y[16]) );
  not_1_47 not_1_component_17 ( .a(a[17]), .y(y[17]) );
  not_1_46 not_1_component_18 ( .a(a[18]), .y(y[18]) );
  not_1_45 not_1_component_19 ( .a(a[19]), .y(y[19]) );
  not_1_44 not_1_component_20 ( .a(a[20]), .y(y[20]) );
  not_1_43 not_1_component_21 ( .a(a[21]), .y(y[21]) );
  not_1_42 not_1_component_22 ( .a(a[22]), .y(y[22]) );
  not_1_41 not_1_component_23 ( .a(a[23]), .y(y[23]) );
  not_1_40 not_1_component_24 ( .a(a[24]), .y(y[24]) );
  not_1_39 not_1_component_25 ( .a(a[25]), .y(y[25]) );
  not_1_38 not_1_component_26 ( .a(a[26]), .y(y[26]) );
  not_1_37 not_1_component_27 ( .a(a[27]), .y(y[27]) );
  not_1_36 not_1_component_28 ( .a(a[28]), .y(y[28]) );
  not_1_35 not_1_component_29 ( .a(a[29]), .y(y[29]) );
  not_1_34 not_1_component_30 ( .a(a[30]), .y(y[30]) );
  not_1_33 not_1_component_31 ( .a(a[31]), .y(y[31]) );
endmodule


module not_1_543 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_542 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_541 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_540 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_539 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_538 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_537 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_536 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_535 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_534 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_533 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_532 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_531 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_530 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_529 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_528 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_527 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_526 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_525 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_524 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_523 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_522 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_521 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_520 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_519 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_518 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_517 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_516 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_515 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_514 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_513 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_512 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_511 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_510 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_509 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_508 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_507 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_506 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_505 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_504 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_503 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_502 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_501 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_500 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_499 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_498 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_497 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_496 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_495 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_494 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_493 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_492 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_491 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_490 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_489 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_488 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_487 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_486 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_485 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_484 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_483 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_482 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_481 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_480 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_479 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_478 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_477 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_476 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_475 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_474 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_473 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_472 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_471 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_470 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_469 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_468 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_467 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_466 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_465 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_464 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_463 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_462 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_461 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_460 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_459 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_458 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_457 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_456 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_455 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_454 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_453 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_452 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_451 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_450 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_449 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_448 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_447 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_446 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_445 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_444 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_443 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_442 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_441 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_440 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_439 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_438 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_437 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_436 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_435 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_434 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_433 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_432 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_431 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_430 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_429 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_428 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_427 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_426 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_425 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_424 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_423 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_422 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_421 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_420 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_419 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_418 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_417 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_416 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_415 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_414 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_413 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_412 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_411 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_410 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_409 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_408 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_407 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_406 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_405 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_404 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_403 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_402 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_401 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_400 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_399 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_398 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_397 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_396 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_395 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_394 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_393 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_392 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_391 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_390 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_389 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_388 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_387 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_386 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_385 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_384 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_383 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_382 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_381 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_380 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_379 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_378 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_377 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_376 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_375 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_374 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_373 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_372 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_371 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_370 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_369 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_368 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_367 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_366 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_365 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_364 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_363 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_362 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_361 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_360 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_359 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_358 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_357 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_356 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_355 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_354 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_353 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_352 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_351 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_350 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_349 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_348 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_347 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_346 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_345 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_344 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_343 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_342 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_341 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_340 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_339 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_338 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_337 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_336 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_335 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_334 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_333 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_332 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_331 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_330 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_329 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_328 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_327 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_326 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_325 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_324 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_323 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_322 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_321 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_320 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_319 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_318 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_317 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_316 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_315 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_314 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_313 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_312 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_311 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_310 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_309 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_308 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_307 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_306 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_305 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_304 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_303 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_302 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_301 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_300 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_299 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_298 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_297 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_296 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_295 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_294 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_293 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_292 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_291 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_290 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_289 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_288 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_287 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_286 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_285 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_284 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_283 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_282 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_281 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_280 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_279 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_278 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_277 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_276 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_275 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_274 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_273 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_272 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_271 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_270 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_269 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_268 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_267 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_266 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_265 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_264 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_263 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_262 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_261 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_260 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_259 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_258 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_257 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_256 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_255 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_254 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_253 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_252 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_251 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_250 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_249 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_248 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_247 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_246 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_245 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_244 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_243 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_242 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_241 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_240 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_239 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_238 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_237 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_236 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_235 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_234 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_233 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_232 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_231 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_230 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_229 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_228 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_227 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_226 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_225 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_224 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_223 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_222 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_221 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_220 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_219 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_218 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_217 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_216 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_215 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_214 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_213 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_212 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_211 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_210 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_209 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_208 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_207 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_206 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_205 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_204 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_203 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_202 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_201 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_200 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_199 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_198 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_197 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_196 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_195 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_194 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_193 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_192 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_191 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_190 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_189 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_188 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_187 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_186 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_185 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_184 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_183 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_182 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_181 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_180 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_179 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_178 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_177 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_176 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_175 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_174 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_173 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_172 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_171 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_170 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_169 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_168 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_167 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_166 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_165 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_164 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_163 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_162 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_161 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_160 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_159 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_158 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_157 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_156 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_155 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_154 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_153 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_152 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_151 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_150 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_149 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_148 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_147 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_146 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_145 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_144 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_143 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_142 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_141 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_140 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_139 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_138 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_137 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_136 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_135 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_134 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_133 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_132 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_131 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_130 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_129 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_128 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_127 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_126 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_125 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_124 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_123 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_122 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_121 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_120 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_119 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_118 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_117 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_116 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_115 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_114 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_113 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_112 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_111 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_110 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_109 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_108 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_107 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_106 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_105 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_104 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_103 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_102 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_101 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_100 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_99 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_98 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_97 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_96 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_95 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_94 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_93 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_92 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_91 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_90 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_89 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_88 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_87 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_86 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_85 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_84 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_83 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_82 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_81 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_80 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_79 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_78 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_77 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_76 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_75 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_74 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_73 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_72 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_71 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_70 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_69 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_68 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_67 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_66 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_65 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_64 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_63 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_62 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_61 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_60 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_59 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_58 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_57 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_56 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_55 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_54 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_53 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_52 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_51 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_50 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_49 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_48 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_47 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_46 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_45 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_44 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_43 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_42 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_41 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_40 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_39 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_38 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_37 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_36 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_35 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_34 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_33 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_32 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_31 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_30 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_29 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_28 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_27 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_26 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_25 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_24 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_23 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_22 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_21 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_20 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_19 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_18 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_17 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_16 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_15 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_14 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_13 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_12 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_11 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_10 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_9 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_8 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_7 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_6 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_5 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_4 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_3 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_2 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module not_1_1 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module or_2_675 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_674 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_673 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_672 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_671 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_670 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_669 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_668 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_667 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_666 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_665 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_664 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_663 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_662 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_661 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_660 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_659 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_658 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_657 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_656 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_655 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_654 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_653 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_652 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_651 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_650 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_649 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_648 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_647 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_646 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_645 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_644 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_643 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_642 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_641 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_640 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_639 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_638 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_637 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_636 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_635 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_634 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_633 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_632 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_631 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_630 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_629 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_628 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_627 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_626 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_625 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_624 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_623 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_622 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_621 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_620 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_619 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_618 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_617 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_616 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_615 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_614 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_613 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_612 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_611 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_610 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_609 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_608 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_607 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_606 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_605 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_604 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_603 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_602 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_601 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_600 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_599 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_598 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_597 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_596 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_595 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_594 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_593 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_592 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_591 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_590 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_589 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_588 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_587 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_586 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_585 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_584 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_583 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_582 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_581 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_580 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_579 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_578 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_577 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_576 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_575 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_574 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_573 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_572 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_571 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_570 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_569 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_568 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_567 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_566 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_565 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_564 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_563 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_562 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_561 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_560 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_559 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_558 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_557 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_556 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_555 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_554 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_553 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_552 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_551 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_550 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_549 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_548 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_547 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_546 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_545 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_544 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_543 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_542 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_541 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_540 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_539 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_538 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_537 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_536 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_535 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_534 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_533 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_532 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_531 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_530 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_529 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_528 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_527 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_526 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_525 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_524 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_523 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_522 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_521 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_520 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_519 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_518 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_517 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_516 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_515 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_514 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_513 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_512 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_511 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_510 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_509 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_508 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_507 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_506 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_505 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_504 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_503 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_502 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_501 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_500 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_499 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_498 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_497 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_496 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_495 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_494 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_493 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_492 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_491 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_490 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_489 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_488 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_487 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_486 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_485 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_484 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_483 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_482 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_481 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_480 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_479 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_478 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_477 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_476 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_475 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_474 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_473 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_472 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_471 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_470 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_469 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_468 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_467 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_466 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_465 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_464 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_463 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_462 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_461 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_460 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_459 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_458 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_457 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_456 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_455 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_454 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_453 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_452 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_451 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_450 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_449 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_448 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_447 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_446 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_445 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_444 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_443 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_442 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_441 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_440 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_439 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_438 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_437 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_436 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_435 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_434 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_433 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_432 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_431 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_430 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_429 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_428 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_427 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_426 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_425 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_424 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_423 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_422 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_421 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_420 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_419 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_418 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_417 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_416 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_415 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_414 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_413 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_412 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_411 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_410 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_409 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_408 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_407 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_406 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_405 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_404 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_403 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_402 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_401 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_400 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_399 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_398 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_397 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_396 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_395 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_394 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_393 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_392 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_391 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_390 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_389 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_388 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_387 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_386 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_385 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_384 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_383 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_382 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_381 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_380 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_379 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_378 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_377 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_376 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_375 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_374 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_373 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_372 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_371 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_370 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_369 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_368 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_367 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_366 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_365 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_364 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_363 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_362 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_361 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_360 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_359 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_358 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_357 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_356 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_355 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_354 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_353 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_352 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_351 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_350 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_349 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_348 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_347 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_346 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_345 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_344 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_343 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_342 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_341 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_340 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_339 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_338 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_337 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_336 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_335 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_334 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_333 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_332 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_331 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_330 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_329 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_328 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_327 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_326 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_325 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_324 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_323 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_322 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_321 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_320 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_319 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_318 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_317 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_316 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_315 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_314 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_313 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_312 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_311 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_310 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_309 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_308 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_307 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_306 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_305 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_304 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_303 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_302 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_301 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_300 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_299 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_298 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_297 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_296 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_295 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_294 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_293 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_292 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_291 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_290 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_289 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_288 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_287 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_286 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_285 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_284 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_283 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_282 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_281 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_280 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_279 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_278 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_277 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_276 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_275 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_274 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_273 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_272 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_271 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_270 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_269 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_268 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_267 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_266 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_265 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_264 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_263 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_262 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_261 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_260 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_259 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_258 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_257 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_256 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_255 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_254 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_253 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_252 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_251 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_250 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_249 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_248 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_247 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_246 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_245 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_244 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_243 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_242 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_241 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_240 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_239 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_238 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_237 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_236 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_235 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_234 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_233 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_232 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_231 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_230 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_229 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_228 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_227 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_226 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_225 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_224 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_223 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_222 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_221 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_220 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_219 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_218 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_217 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_216 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_215 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_214 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_213 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_212 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_211 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_210 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_209 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_208 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_207 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_206 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_205 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_204 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_203 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_202 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_201 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_200 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_199 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_198 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_197 ( a, b, y );
  input a, b;
  output y;

  tri   y;

  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_196 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_195 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_194 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_193 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_192 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_191 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_190 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_189 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_188 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_187 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_186 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_185 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_184 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_183 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_182 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_181 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_180 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_179 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_178 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_177 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_176 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_175 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_174 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_173 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_172 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_171 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_170 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_169 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_168 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_167 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_166 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_165 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_164 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_163 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_162 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_161 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_160 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_159 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_158 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_157 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_156 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_155 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_154 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_153 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_152 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_151 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_150 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_149 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_148 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_147 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_146 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_145 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_144 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_143 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_142 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_141 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_140 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_139 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_138 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_137 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_136 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_135 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_134 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_133 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_132 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_131 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_130 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_129 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_128 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_127 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_126 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_125 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_124 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_123 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_122 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_121 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_120 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_119 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_118 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_117 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_116 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_115 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_114 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_113 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_112 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_111 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_110 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_109 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_108 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_107 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_106 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_105 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_104 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_103 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_102 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_101 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_100 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_99 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_98 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_97 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_96 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_95 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_94 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_93 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_92 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_91 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_90 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_89 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_88 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_87 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_86 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_85 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_84 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_83 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_82 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_81 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_80 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_79 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_78 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_77 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_76 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_75 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_74 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_73 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_72 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_71 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_70 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_69 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_68 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_67 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_66 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_65 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_64 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_63 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_62 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_61 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_60 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_59 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_58 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_57 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_56 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_55 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_54 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_53 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_52 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_51 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_50 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_49 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_48 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_47 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_46 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_45 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_44 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_43 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_42 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_41 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_40 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_39 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_38 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_37 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_36 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_35 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_34 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_33 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_32 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_31 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_30 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_29 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_28 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_27 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_26 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_25 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_24 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_23 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_22 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_21 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_20 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_19 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_18 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_17 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_16 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_15 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_14 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_13 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_12 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_11 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_10 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_9 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_8 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_7 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_6 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_5 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_4 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_3 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_2 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module or_2_1 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module mux21_479 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_543 inv ( .a(s), .y(sa) );
  and_2_1309 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1308 and2 ( .a(b), .b(s), .y(y2) );
  or_2_643 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_478 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_542 inv ( .a(s), .y(sa) );
  and_2_1307 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1306 and2 ( .a(b), .b(s), .y(y2) );
  or_2_642 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_477 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_541 inv ( .a(s), .y(sa) );
  and_2_1305 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1304 and2 ( .a(b), .b(s), .y(y2) );
  or_2_641 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_476 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_540 inv ( .a(s), .y(sa) );
  and_2_1303 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1302 and2 ( .a(b), .b(s), .y(y2) );
  or_2_640 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_475 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_539 inv ( .a(s), .y(sa) );
  and_2_1301 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1300 and2 ( .a(b), .b(s), .y(y2) );
  or_2_639 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_474 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_538 inv ( .a(s), .y(sa) );
  and_2_1299 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1298 and2 ( .a(b), .b(s), .y(y2) );
  or_2_638 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_473 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_537 inv ( .a(s), .y(sa) );
  and_2_1297 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1296 and2 ( .a(b), .b(s), .y(y2) );
  or_2_637 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_472 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_536 inv ( .a(s), .y(sa) );
  and_2_1295 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1294 and2 ( .a(b), .b(s), .y(y2) );
  or_2_636 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_471 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_535 inv ( .a(s), .y(sa) );
  and_2_1293 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1292 and2 ( .a(b), .b(s), .y(y2) );
  or_2_635 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_470 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_534 inv ( .a(s), .y(sa) );
  and_2_1291 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1290 and2 ( .a(b), .b(s), .y(y2) );
  or_2_634 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_469 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_533 inv ( .a(s), .y(sa) );
  and_2_1289 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1288 and2 ( .a(b), .b(s), .y(y2) );
  or_2_633 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_468 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_532 inv ( .a(s), .y(sa) );
  and_2_1287 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1286 and2 ( .a(b), .b(s), .y(y2) );
  or_2_632 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_467 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_531 inv ( .a(s), .y(sa) );
  and_2_1285 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1284 and2 ( .a(b), .b(s), .y(y2) );
  or_2_631 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_466 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_530 inv ( .a(s), .y(sa) );
  and_2_1283 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1282 and2 ( .a(b), .b(s), .y(y2) );
  or_2_630 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_465 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_529 inv ( .a(s), .y(sa) );
  and_2_1281 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1280 and2 ( .a(b), .b(s), .y(y2) );
  or_2_629 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_464 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_528 inv ( .a(s), .y(sa) );
  and_2_1279 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1278 and2 ( .a(b), .b(s), .y(y2) );
  or_2_628 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_463 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_527 inv ( .a(s), .y(sa) );
  and_2_1277 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1276 and2 ( .a(b), .b(s), .y(y2) );
  or_2_627 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_462 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_526 inv ( .a(s), .y(sa) );
  and_2_1275 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1274 and2 ( .a(b), .b(s), .y(y2) );
  or_2_626 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_461 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_525 inv ( .a(s), .y(sa) );
  and_2_1273 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1272 and2 ( .a(b), .b(s), .y(y2) );
  or_2_625 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_460 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_524 inv ( .a(s), .y(sa) );
  and_2_1271 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1270 and2 ( .a(b), .b(s), .y(y2) );
  or_2_624 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_459 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_523 inv ( .a(s), .y(sa) );
  and_2_1269 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1268 and2 ( .a(b), .b(s), .y(y2) );
  or_2_623 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_458 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_522 inv ( .a(s), .y(sa) );
  and_2_1267 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1266 and2 ( .a(b), .b(s), .y(y2) );
  or_2_622 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_457 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_521 inv ( .a(s), .y(sa) );
  and_2_1265 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1264 and2 ( .a(b), .b(s), .y(y2) );
  or_2_621 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_456 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_520 inv ( .a(s), .y(sa) );
  and_2_1263 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1262 and2 ( .a(b), .b(s), .y(y2) );
  or_2_620 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_455 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_519 inv ( .a(s), .y(sa) );
  and_2_1261 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1260 and2 ( .a(b), .b(s), .y(y2) );
  or_2_619 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_454 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_518 inv ( .a(s), .y(sa) );
  and_2_1259 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1258 and2 ( .a(b), .b(s), .y(y2) );
  or_2_618 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_453 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_517 inv ( .a(s), .y(sa) );
  and_2_1257 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1256 and2 ( .a(b), .b(s), .y(y2) );
  or_2_617 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_452 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_516 inv ( .a(s), .y(sa) );
  and_2_1255 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1254 and2 ( .a(b), .b(s), .y(y2) );
  or_2_616 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_451 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_515 inv ( .a(s), .y(sa) );
  and_2_1253 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1252 and2 ( .a(b), .b(s), .y(y2) );
  or_2_615 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_450 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_514 inv ( .a(s), .y(sa) );
  and_2_1251 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1250 and2 ( .a(b), .b(s), .y(y2) );
  or_2_614 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_449 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_513 inv ( .a(s), .y(sa) );
  and_2_1249 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1248 and2 ( .a(b), .b(s), .y(y2) );
  or_2_613 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_448 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_512 inv ( .a(s), .y(sa) );
  and_2_1247 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1246 and2 ( .a(b), .b(s), .y(y2) );
  or_2_612 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_447 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_511 inv ( .a(s), .y(sa) );
  and_2_1245 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1244 and2 ( .a(b), .b(s), .y(y2) );
  or_2_611 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_446 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_510 inv ( .a(s), .y(sa) );
  and_2_1243 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1242 and2 ( .a(b), .b(s), .y(y2) );
  or_2_610 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_445 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_509 inv ( .a(s), .y(sa) );
  and_2_1241 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1240 and2 ( .a(b), .b(s), .y(y2) );
  or_2_609 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_444 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_508 inv ( .a(s), .y(sa) );
  and_2_1239 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1238 and2 ( .a(b), .b(s), .y(y2) );
  or_2_608 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_443 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_507 inv ( .a(s), .y(sa) );
  and_2_1237 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1236 and2 ( .a(b), .b(s), .y(y2) );
  or_2_607 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_442 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_506 inv ( .a(s), .y(sa) );
  and_2_1235 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1234 and2 ( .a(b), .b(s), .y(y2) );
  or_2_606 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_441 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_505 inv ( .a(s), .y(sa) );
  and_2_1233 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1232 and2 ( .a(b), .b(s), .y(y2) );
  or_2_605 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_440 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_504 inv ( .a(s), .y(sa) );
  and_2_1231 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1230 and2 ( .a(b), .b(s), .y(y2) );
  or_2_604 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_439 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_503 inv ( .a(s), .y(sa) );
  and_2_1229 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1228 and2 ( .a(b), .b(s), .y(y2) );
  or_2_603 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_438 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_502 inv ( .a(s), .y(sa) );
  and_2_1227 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1226 and2 ( .a(b), .b(s), .y(y2) );
  or_2_602 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_437 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_501 inv ( .a(s), .y(sa) );
  and_2_1225 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1224 and2 ( .a(b), .b(s), .y(y2) );
  or_2_601 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_436 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_500 inv ( .a(s), .y(sa) );
  and_2_1223 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1222 and2 ( .a(b), .b(s), .y(y2) );
  or_2_600 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_435 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_499 inv ( .a(s), .y(sa) );
  and_2_1221 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1220 and2 ( .a(b), .b(s), .y(y2) );
  or_2_599 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_434 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_498 inv ( .a(s), .y(sa) );
  and_2_1219 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1218 and2 ( .a(b), .b(s), .y(y2) );
  or_2_598 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_433 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_497 inv ( .a(s), .y(sa) );
  and_2_1217 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1216 and2 ( .a(b), .b(s), .y(y2) );
  or_2_597 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_432 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_496 inv ( .a(s), .y(sa) );
  and_2_1215 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1214 and2 ( .a(b), .b(s), .y(y2) );
  or_2_596 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_431 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_495 inv ( .a(s), .y(sa) );
  and_2_1213 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1212 and2 ( .a(b), .b(s), .y(y2) );
  or_2_595 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_430 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_494 inv ( .a(s), .y(sa) );
  and_2_1211 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1210 and2 ( .a(b), .b(s), .y(y2) );
  or_2_594 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_429 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_493 inv ( .a(s), .y(sa) );
  and_2_1209 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1208 and2 ( .a(b), .b(s), .y(y2) );
  or_2_593 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_428 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_492 inv ( .a(s), .y(sa) );
  and_2_1207 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1206 and2 ( .a(b), .b(s), .y(y2) );
  or_2_592 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_427 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_491 inv ( .a(s), .y(sa) );
  and_2_1205 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1204 and2 ( .a(b), .b(s), .y(y2) );
  or_2_591 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_426 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_490 inv ( .a(s), .y(sa) );
  and_2_1203 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1202 and2 ( .a(b), .b(s), .y(y2) );
  or_2_590 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_425 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_489 inv ( .a(s), .y(sa) );
  and_2_1201 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1200 and2 ( .a(b), .b(s), .y(y2) );
  or_2_589 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_424 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_488 inv ( .a(s), .y(sa) );
  and_2_1199 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1198 and2 ( .a(b), .b(s), .y(y2) );
  or_2_588 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_423 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_487 inv ( .a(s), .y(sa) );
  and_2_1197 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1196 and2 ( .a(b), .b(s), .y(y2) );
  or_2_587 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_422 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_486 inv ( .a(s), .y(sa) );
  and_2_1195 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1194 and2 ( .a(b), .b(s), .y(y2) );
  or_2_586 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_421 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_485 inv ( .a(s), .y(sa) );
  and_2_1193 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1192 and2 ( .a(b), .b(s), .y(y2) );
  or_2_585 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_420 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_484 inv ( .a(s), .y(sa) );
  and_2_1191 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1190 and2 ( .a(b), .b(s), .y(y2) );
  or_2_584 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_419 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_483 inv ( .a(s), .y(sa) );
  and_2_1189 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1188 and2 ( .a(b), .b(s), .y(y2) );
  or_2_583 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_418 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_482 inv ( .a(s), .y(sa) );
  and_2_1187 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1186 and2 ( .a(b), .b(s), .y(y2) );
  or_2_582 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_417 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_481 inv ( .a(s), .y(sa) );
  and_2_1185 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1184 and2 ( .a(b), .b(s), .y(y2) );
  or_2_581 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_416 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_480 inv ( .a(s), .y(sa) );
  and_2_1183 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1182 and2 ( .a(b), .b(s), .y(y2) );
  or_2_580 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_415 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_479 inv ( .a(s), .y(sa) );
  and_2_1181 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1180 and2 ( .a(b), .b(s), .y(y2) );
  or_2_579 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_414 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_478 inv ( .a(s), .y(sa) );
  and_2_1179 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1178 and2 ( .a(b), .b(s), .y(y2) );
  or_2_578 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_413 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_477 inv ( .a(s), .y(sa) );
  and_2_1177 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1176 and2 ( .a(b), .b(s), .y(y2) );
  or_2_577 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_412 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_476 inv ( .a(s), .y(sa) );
  and_2_1175 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1174 and2 ( .a(b), .b(s), .y(y2) );
  or_2_576 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_411 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_475 inv ( .a(s), .y(sa) );
  and_2_1173 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1172 and2 ( .a(b), .b(s), .y(y2) );
  or_2_575 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_410 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_474 inv ( .a(s), .y(sa) );
  and_2_1171 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1170 and2 ( .a(b), .b(s), .y(y2) );
  or_2_574 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_409 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_473 inv ( .a(s), .y(sa) );
  and_2_1169 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1168 and2 ( .a(b), .b(s), .y(y2) );
  or_2_573 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_408 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_472 inv ( .a(s), .y(sa) );
  and_2_1167 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1166 and2 ( .a(b), .b(s), .y(y2) );
  or_2_572 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_407 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_471 inv ( .a(s), .y(sa) );
  and_2_1165 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1164 and2 ( .a(b), .b(s), .y(y2) );
  or_2_571 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_406 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_470 inv ( .a(s), .y(sa) );
  and_2_1163 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1162 and2 ( .a(b), .b(s), .y(y2) );
  or_2_570 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_405 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_469 inv ( .a(s), .y(sa) );
  and_2_1161 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1160 and2 ( .a(b), .b(s), .y(y2) );
  or_2_569 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_404 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_468 inv ( .a(s), .y(sa) );
  and_2_1159 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1158 and2 ( .a(b), .b(s), .y(y2) );
  or_2_568 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_403 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_467 inv ( .a(s), .y(sa) );
  and_2_1157 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1156 and2 ( .a(b), .b(s), .y(y2) );
  or_2_567 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_402 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_466 inv ( .a(s), .y(sa) );
  and_2_1155 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1154 and2 ( .a(b), .b(s), .y(y2) );
  or_2_566 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_401 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_465 inv ( .a(s), .y(sa) );
  and_2_1153 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1152 and2 ( .a(b), .b(s), .y(y2) );
  or_2_565 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_400 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_464 inv ( .a(s), .y(sa) );
  and_2_1151 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1150 and2 ( .a(b), .b(s), .y(y2) );
  or_2_564 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_399 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_463 inv ( .a(s), .y(sa) );
  and_2_1149 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1148 and2 ( .a(b), .b(s), .y(y2) );
  or_2_563 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_398 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_462 inv ( .a(s), .y(sa) );
  and_2_1147 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1146 and2 ( .a(b), .b(s), .y(y2) );
  or_2_562 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_397 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_461 inv ( .a(s), .y(sa) );
  and_2_1145 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1144 and2 ( .a(b), .b(s), .y(y2) );
  or_2_561 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_396 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_460 inv ( .a(s), .y(sa) );
  and_2_1143 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1142 and2 ( .a(b), .b(s), .y(y2) );
  or_2_560 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_395 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_459 inv ( .a(s), .y(sa) );
  and_2_1141 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1140 and2 ( .a(b), .b(s), .y(y2) );
  or_2_559 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_394 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_458 inv ( .a(s), .y(sa) );
  and_2_1139 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1138 and2 ( .a(b), .b(s), .y(y2) );
  or_2_558 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_393 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_457 inv ( .a(s), .y(sa) );
  and_2_1137 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1136 and2 ( .a(b), .b(s), .y(y2) );
  or_2_557 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_392 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_456 inv ( .a(s), .y(sa) );
  and_2_1135 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1134 and2 ( .a(b), .b(s), .y(y2) );
  or_2_556 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_391 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_455 inv ( .a(s), .y(sa) );
  and_2_1133 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1132 and2 ( .a(b), .b(s), .y(y2) );
  or_2_555 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_390 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_454 inv ( .a(s), .y(sa) );
  and_2_1131 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1130 and2 ( .a(b), .b(s), .y(y2) );
  or_2_554 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_389 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_453 inv ( .a(s), .y(sa) );
  and_2_1129 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1128 and2 ( .a(b), .b(s), .y(y2) );
  or_2_553 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_388 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_452 inv ( .a(s), .y(sa) );
  and_2_1127 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1126 and2 ( .a(b), .b(s), .y(y2) );
  or_2_552 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_387 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_451 inv ( .a(s), .y(sa) );
  and_2_1125 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1124 and2 ( .a(b), .b(s), .y(y2) );
  or_2_551 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_386 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_450 inv ( .a(s), .y(sa) );
  and_2_1123 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1122 and2 ( .a(b), .b(s), .y(y2) );
  or_2_550 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_385 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_449 inv ( .a(s), .y(sa) );
  and_2_1121 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1120 and2 ( .a(b), .b(s), .y(y2) );
  or_2_549 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_384 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_448 inv ( .a(s), .y(sa) );
  and_2_1119 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1118 and2 ( .a(b), .b(s), .y(y2) );
  or_2_548 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_383 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_447 inv ( .a(s), .y(sa) );
  and_2_1117 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1116 and2 ( .a(b), .b(s), .y(y2) );
  or_2_547 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_382 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_446 inv ( .a(s), .y(sa) );
  and_2_1115 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1114 and2 ( .a(b), .b(s), .y(y2) );
  or_2_546 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_381 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_445 inv ( .a(s), .y(sa) );
  and_2_1113 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1112 and2 ( .a(b), .b(s), .y(y2) );
  or_2_545 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_380 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_444 inv ( .a(s), .y(sa) );
  and_2_1111 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1110 and2 ( .a(b), .b(s), .y(y2) );
  or_2_544 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_379 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_443 inv ( .a(s), .y(sa) );
  and_2_1109 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1108 and2 ( .a(b), .b(s), .y(y2) );
  or_2_543 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_378 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_442 inv ( .a(s), .y(sa) );
  and_2_1107 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1106 and2 ( .a(b), .b(s), .y(y2) );
  or_2_542 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_377 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_441 inv ( .a(s), .y(sa) );
  and_2_1105 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1104 and2 ( .a(b), .b(s), .y(y2) );
  or_2_541 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_376 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_440 inv ( .a(s), .y(sa) );
  and_2_1103 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1102 and2 ( .a(b), .b(s), .y(y2) );
  or_2_540 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_375 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_439 inv ( .a(s), .y(sa) );
  and_2_1101 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1100 and2 ( .a(b), .b(s), .y(y2) );
  or_2_539 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_374 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_438 inv ( .a(s), .y(sa) );
  and_2_1099 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1098 and2 ( .a(b), .b(s), .y(y2) );
  or_2_538 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_373 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_437 inv ( .a(s), .y(sa) );
  and_2_1097 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1096 and2 ( .a(b), .b(s), .y(y2) );
  or_2_537 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_372 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_436 inv ( .a(s), .y(sa) );
  and_2_1095 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1094 and2 ( .a(b), .b(s), .y(y2) );
  or_2_536 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_371 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_435 inv ( .a(s), .y(sa) );
  and_2_1093 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1092 and2 ( .a(b), .b(s), .y(y2) );
  or_2_535 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_370 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_434 inv ( .a(s), .y(sa) );
  and_2_1091 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1090 and2 ( .a(b), .b(s), .y(y2) );
  or_2_534 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_369 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_433 inv ( .a(s), .y(sa) );
  and_2_1089 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1088 and2 ( .a(b), .b(s), .y(y2) );
  or_2_533 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_368 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_432 inv ( .a(s), .y(sa) );
  and_2_1087 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1086 and2 ( .a(b), .b(s), .y(y2) );
  or_2_532 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_367 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_431 inv ( .a(s), .y(sa) );
  and_2_1085 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1084 and2 ( .a(b), .b(s), .y(y2) );
  or_2_531 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_366 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_430 inv ( .a(s), .y(sa) );
  and_2_1083 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1082 and2 ( .a(b), .b(s), .y(y2) );
  or_2_530 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_365 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_429 inv ( .a(s), .y(sa) );
  and_2_1081 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1080 and2 ( .a(b), .b(s), .y(y2) );
  or_2_529 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_364 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_428 inv ( .a(s), .y(sa) );
  and_2_1079 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1078 and2 ( .a(b), .b(s), .y(y2) );
  or_2_528 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_363 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_427 inv ( .a(s), .y(sa) );
  and_2_1077 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1076 and2 ( .a(b), .b(s), .y(y2) );
  or_2_527 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_362 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_426 inv ( .a(s), .y(sa) );
  and_2_1075 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1074 and2 ( .a(b), .b(s), .y(y2) );
  or_2_526 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_361 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_425 inv ( .a(s), .y(sa) );
  and_2_1073 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1072 and2 ( .a(b), .b(s), .y(y2) );
  or_2_525 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_360 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_424 inv ( .a(s), .y(sa) );
  and_2_1071 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1070 and2 ( .a(b), .b(s), .y(y2) );
  or_2_524 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_359 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_423 inv ( .a(s), .y(sa) );
  and_2_1069 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1068 and2 ( .a(b), .b(s), .y(y2) );
  or_2_523 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_358 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_422 inv ( .a(s), .y(sa) );
  and_2_1067 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1066 and2 ( .a(b), .b(s), .y(y2) );
  or_2_522 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_357 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_421 inv ( .a(s), .y(sa) );
  and_2_1065 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1064 and2 ( .a(b), .b(s), .y(y2) );
  or_2_521 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_356 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_420 inv ( .a(s), .y(sa) );
  and_2_1063 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1062 and2 ( .a(b), .b(s), .y(y2) );
  or_2_520 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_355 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_419 inv ( .a(s), .y(sa) );
  and_2_1061 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1060 and2 ( .a(b), .b(s), .y(y2) );
  or_2_519 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_354 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_418 inv ( .a(s), .y(sa) );
  and_2_1059 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1058 and2 ( .a(b), .b(s), .y(y2) );
  or_2_518 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_353 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_417 inv ( .a(s), .y(sa) );
  and_2_1057 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1056 and2 ( .a(b), .b(s), .y(y2) );
  or_2_517 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_352 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_384 inv ( .a(s), .y(sa) );
  and_2_1055 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1054 and2 ( .a(b), .b(s), .y(y2) );
  or_2_516 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_351 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_383 inv ( .a(s), .y(sa) );
  and_2_1053 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1052 and2 ( .a(b), .b(s), .y(y2) );
  or_2_515 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_350 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_382 inv ( .a(s), .y(sa) );
  and_2_1051 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1050 and2 ( .a(b), .b(s), .y(y2) );
  or_2_514 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_349 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_381 inv ( .a(s), .y(sa) );
  and_2_1049 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1048 and2 ( .a(b), .b(s), .y(y2) );
  or_2_513 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_348 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_380 inv ( .a(s), .y(sa) );
  and_2_1047 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1046 and2 ( .a(b), .b(s), .y(y2) );
  or_2_512 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_347 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_379 inv ( .a(s), .y(sa) );
  and_2_1045 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1044 and2 ( .a(b), .b(s), .y(y2) );
  or_2_511 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_346 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_378 inv ( .a(s), .y(sa) );
  and_2_1043 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1042 and2 ( .a(b), .b(s), .y(y2) );
  or_2_510 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_345 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_377 inv ( .a(s), .y(sa) );
  and_2_1041 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1040 and2 ( .a(b), .b(s), .y(y2) );
  or_2_509 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_344 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_376 inv ( .a(s), .y(sa) );
  and_2_1039 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1038 and2 ( .a(b), .b(s), .y(y2) );
  or_2_508 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_343 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_375 inv ( .a(s), .y(sa) );
  and_2_1037 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1036 and2 ( .a(b), .b(s), .y(y2) );
  or_2_507 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_342 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_374 inv ( .a(s), .y(sa) );
  and_2_1035 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1034 and2 ( .a(b), .b(s), .y(y2) );
  or_2_506 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_341 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_373 inv ( .a(s), .y(sa) );
  and_2_1033 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1032 and2 ( .a(b), .b(s), .y(y2) );
  or_2_505 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_340 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_372 inv ( .a(s), .y(sa) );
  and_2_1031 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1030 and2 ( .a(b), .b(s), .y(y2) );
  or_2_504 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_339 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_371 inv ( .a(s), .y(sa) );
  and_2_1029 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1028 and2 ( .a(b), .b(s), .y(y2) );
  or_2_503 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_338 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_370 inv ( .a(s), .y(sa) );
  and_2_1027 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1026 and2 ( .a(b), .b(s), .y(y2) );
  or_2_502 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_337 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_369 inv ( .a(s), .y(sa) );
  and_2_1025 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1024 and2 ( .a(b), .b(s), .y(y2) );
  or_2_501 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_336 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_368 inv ( .a(s), .y(sa) );
  and_2_1023 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1022 and2 ( .a(b), .b(s), .y(y2) );
  or_2_500 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_335 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_367 inv ( .a(s), .y(sa) );
  and_2_1021 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1020 and2 ( .a(b), .b(s), .y(y2) );
  or_2_499 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_334 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_366 inv ( .a(s), .y(sa) );
  and_2_1019 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1018 and2 ( .a(b), .b(s), .y(y2) );
  or_2_498 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_333 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_365 inv ( .a(s), .y(sa) );
  and_2_1017 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1016 and2 ( .a(b), .b(s), .y(y2) );
  or_2_497 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_332 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_364 inv ( .a(s), .y(sa) );
  and_2_1015 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1014 and2 ( .a(b), .b(s), .y(y2) );
  or_2_496 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_331 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_363 inv ( .a(s), .y(sa) );
  and_2_1013 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1012 and2 ( .a(b), .b(s), .y(y2) );
  or_2_495 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_330 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_362 inv ( .a(s), .y(sa) );
  and_2_1011 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1010 and2 ( .a(b), .b(s), .y(y2) );
  or_2_494 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_329 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_361 inv ( .a(s), .y(sa) );
  and_2_1009 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1008 and2 ( .a(b), .b(s), .y(y2) );
  or_2_493 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_328 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_360 inv ( .a(s), .y(sa) );
  and_2_1007 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1006 and2 ( .a(b), .b(s), .y(y2) );
  or_2_492 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_327 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_359 inv ( .a(s), .y(sa) );
  and_2_1005 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1004 and2 ( .a(b), .b(s), .y(y2) );
  or_2_491 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_326 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_358 inv ( .a(s), .y(sa) );
  and_2_1003 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1002 and2 ( .a(b), .b(s), .y(y2) );
  or_2_490 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_325 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_357 inv ( .a(s), .y(sa) );
  and_2_1001 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1000 and2 ( .a(b), .b(s), .y(y2) );
  or_2_489 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_324 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_356 inv ( .a(s), .y(sa) );
  and_2_999 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_998 and2 ( .a(b), .b(s), .y(y2) );
  or_2_488 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_323 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_355 inv ( .a(s), .y(sa) );
  and_2_997 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_996 and2 ( .a(b), .b(s), .y(y2) );
  or_2_487 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_322 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_354 inv ( .a(s), .y(sa) );
  and_2_995 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_994 and2 ( .a(b), .b(s), .y(y2) );
  or_2_486 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_321 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_353 inv ( .a(s), .y(sa) );
  and_2_993 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_992 and2 ( .a(b), .b(s), .y(y2) );
  or_2_485 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_320 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_352 inv ( .a(s), .y(sa) );
  and_2_991 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_990 and2 ( .a(b), .b(s), .y(y2) );
  or_2_484 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_319 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_351 inv ( .a(s), .y(sa) );
  and_2_989 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_988 and2 ( .a(b), .b(s), .y(y2) );
  or_2_483 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_318 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_350 inv ( .a(s), .y(sa) );
  and_2_987 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_986 and2 ( .a(b), .b(s), .y(y2) );
  or_2_482 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_317 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_349 inv ( .a(s), .y(sa) );
  and_2_985 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_984 and2 ( .a(b), .b(s), .y(y2) );
  or_2_481 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_316 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_348 inv ( .a(s), .y(sa) );
  and_2_983 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_982 and2 ( .a(b), .b(s), .y(y2) );
  or_2_480 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_315 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_347 inv ( .a(s), .y(sa) );
  and_2_981 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_980 and2 ( .a(b), .b(s), .y(y2) );
  or_2_479 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_314 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_346 inv ( .a(s), .y(sa) );
  and_2_979 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_978 and2 ( .a(b), .b(s), .y(y2) );
  or_2_478 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_313 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_345 inv ( .a(s), .y(sa) );
  and_2_977 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_976 and2 ( .a(b), .b(s), .y(y2) );
  or_2_477 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_312 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_344 inv ( .a(s), .y(sa) );
  and_2_975 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_974 and2 ( .a(b), .b(s), .y(y2) );
  or_2_476 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_311 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_343 inv ( .a(s), .y(sa) );
  and_2_973 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_972 and2 ( .a(b), .b(s), .y(y2) );
  or_2_475 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_310 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_342 inv ( .a(s), .y(sa) );
  and_2_971 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_970 and2 ( .a(b), .b(s), .y(y2) );
  or_2_474 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_309 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_341 inv ( .a(s), .y(sa) );
  and_2_969 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_968 and2 ( .a(b), .b(s), .y(y2) );
  or_2_473 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_308 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_340 inv ( .a(s), .y(sa) );
  and_2_967 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_966 and2 ( .a(b), .b(s), .y(y2) );
  or_2_472 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_307 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_339 inv ( .a(s), .y(sa) );
  and_2_965 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_964 and2 ( .a(b), .b(s), .y(y2) );
  or_2_471 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_306 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_338 inv ( .a(s), .y(sa) );
  and_2_963 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_962 and2 ( .a(b), .b(s), .y(y2) );
  or_2_470 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_305 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_337 inv ( .a(s), .y(sa) );
  and_2_961 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_960 and2 ( .a(b), .b(s), .y(y2) );
  or_2_469 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_304 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_336 inv ( .a(s), .y(sa) );
  and_2_959 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_958 and2 ( .a(b), .b(s), .y(y2) );
  or_2_468 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_303 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_335 inv ( .a(s), .y(sa) );
  and_2_957 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_956 and2 ( .a(b), .b(s), .y(y2) );
  or_2_467 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_302 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_334 inv ( .a(s), .y(sa) );
  and_2_955 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_954 and2 ( .a(b), .b(s), .y(y2) );
  or_2_466 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_301 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_333 inv ( .a(s), .y(sa) );
  and_2_953 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_952 and2 ( .a(b), .b(s), .y(y2) );
  or_2_465 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_300 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_332 inv ( .a(s), .y(sa) );
  and_2_951 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_950 and2 ( .a(b), .b(s), .y(y2) );
  or_2_464 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_299 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_331 inv ( .a(s), .y(sa) );
  and_2_949 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_948 and2 ( .a(b), .b(s), .y(y2) );
  or_2_463 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_298 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_330 inv ( .a(s), .y(sa) );
  and_2_947 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_946 and2 ( .a(b), .b(s), .y(y2) );
  or_2_462 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_297 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_329 inv ( .a(s), .y(sa) );
  and_2_945 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_944 and2 ( .a(b), .b(s), .y(y2) );
  or_2_461 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_296 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_328 inv ( .a(s), .y(sa) );
  and_2_943 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_942 and2 ( .a(b), .b(s), .y(y2) );
  or_2_460 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_295 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_327 inv ( .a(s), .y(sa) );
  and_2_941 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_940 and2 ( .a(b), .b(s), .y(y2) );
  or_2_459 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_294 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_326 inv ( .a(s), .y(sa) );
  and_2_939 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_938 and2 ( .a(b), .b(s), .y(y2) );
  or_2_458 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_293 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_325 inv ( .a(s), .y(sa) );
  and_2_937 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_936 and2 ( .a(b), .b(s), .y(y2) );
  or_2_457 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_292 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_324 inv ( .a(s), .y(sa) );
  and_2_935 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_934 and2 ( .a(b), .b(s), .y(y2) );
  or_2_456 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_291 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_323 inv ( .a(s), .y(sa) );
  and_2_933 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_932 and2 ( .a(b), .b(s), .y(y2) );
  or_2_455 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_290 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_322 inv ( .a(s), .y(sa) );
  and_2_931 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_930 and2 ( .a(b), .b(s), .y(y2) );
  or_2_454 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_289 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_321 inv ( .a(s), .y(sa) );
  and_2_929 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_928 and2 ( .a(b), .b(s), .y(y2) );
  or_2_453 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_288 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_320 inv ( .a(s), .y(sa) );
  and_2_927 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_926 and2 ( .a(b), .b(s), .y(y2) );
  or_2_452 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_287 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_319 inv ( .a(s), .y(sa) );
  and_2_925 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_924 and2 ( .a(b), .b(s), .y(y2) );
  or_2_451 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_286 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_318 inv ( .a(s), .y(sa) );
  and_2_923 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_922 and2 ( .a(b), .b(s), .y(y2) );
  or_2_450 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_285 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_317 inv ( .a(s), .y(sa) );
  and_2_921 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_920 and2 ( .a(b), .b(s), .y(y2) );
  or_2_449 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_284 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_316 inv ( .a(s), .y(sa) );
  and_2_919 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_918 and2 ( .a(b), .b(s), .y(y2) );
  or_2_448 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_283 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_315 inv ( .a(s), .y(sa) );
  and_2_917 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_916 and2 ( .a(b), .b(s), .y(y2) );
  or_2_447 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_282 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_314 inv ( .a(s), .y(sa) );
  and_2_915 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_914 and2 ( .a(b), .b(s), .y(y2) );
  or_2_446 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_281 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_313 inv ( .a(s), .y(sa) );
  and_2_913 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_912 and2 ( .a(b), .b(s), .y(y2) );
  or_2_445 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_280 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_312 inv ( .a(s), .y(sa) );
  and_2_911 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_910 and2 ( .a(b), .b(s), .y(y2) );
  or_2_444 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_279 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_311 inv ( .a(s), .y(sa) );
  and_2_909 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_908 and2 ( .a(b), .b(s), .y(y2) );
  or_2_443 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_278 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_310 inv ( .a(s), .y(sa) );
  and_2_907 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_906 and2 ( .a(b), .b(s), .y(y2) );
  or_2_442 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_277 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_309 inv ( .a(s), .y(sa) );
  and_2_905 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_904 and2 ( .a(b), .b(s), .y(y2) );
  or_2_441 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_276 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_308 inv ( .a(s), .y(sa) );
  and_2_903 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_902 and2 ( .a(b), .b(s), .y(y2) );
  or_2_440 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_275 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_307 inv ( .a(s), .y(sa) );
  and_2_901 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_900 and2 ( .a(b), .b(s), .y(y2) );
  or_2_439 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_274 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_306 inv ( .a(s), .y(sa) );
  and_2_899 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_898 and2 ( .a(b), .b(s), .y(y2) );
  or_2_438 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_273 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_305 inv ( .a(s), .y(sa) );
  and_2_897 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_896 and2 ( .a(b), .b(s), .y(y2) );
  or_2_437 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_272 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_304 inv ( .a(s), .y(sa) );
  and_2_895 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_894 and2 ( .a(b), .b(s), .y(y2) );
  or_2_436 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_271 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_303 inv ( .a(s), .y(sa) );
  and_2_893 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_892 and2 ( .a(b), .b(s), .y(y2) );
  or_2_435 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_270 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_302 inv ( .a(s), .y(sa) );
  and_2_891 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_890 and2 ( .a(b), .b(s), .y(y2) );
  or_2_434 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_269 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_301 inv ( .a(s), .y(sa) );
  and_2_889 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_888 and2 ( .a(b), .b(s), .y(y2) );
  or_2_433 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_268 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_300 inv ( .a(s), .y(sa) );
  and_2_887 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_886 and2 ( .a(b), .b(s), .y(y2) );
  or_2_432 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_267 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_299 inv ( .a(s), .y(sa) );
  and_2_885 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_884 and2 ( .a(b), .b(s), .y(y2) );
  or_2_431 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_266 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_298 inv ( .a(s), .y(sa) );
  and_2_883 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_882 and2 ( .a(b), .b(s), .y(y2) );
  or_2_430 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_265 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_297 inv ( .a(s), .y(sa) );
  and_2_881 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_880 and2 ( .a(b), .b(s), .y(y2) );
  or_2_429 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_264 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_296 inv ( .a(s), .y(sa) );
  and_2_879 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_878 and2 ( .a(b), .b(s), .y(y2) );
  or_2_428 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_263 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_295 inv ( .a(s), .y(sa) );
  and_2_877 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_876 and2 ( .a(b), .b(s), .y(y2) );
  or_2_427 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_262 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_294 inv ( .a(s), .y(sa) );
  and_2_875 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_874 and2 ( .a(b), .b(s), .y(y2) );
  or_2_426 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_261 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_293 inv ( .a(s), .y(sa) );
  and_2_873 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_872 and2 ( .a(b), .b(s), .y(y2) );
  or_2_425 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_260 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_292 inv ( .a(s), .y(sa) );
  and_2_871 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_870 and2 ( .a(b), .b(s), .y(y2) );
  or_2_424 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_259 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_291 inv ( .a(s), .y(sa) );
  and_2_869 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_868 and2 ( .a(b), .b(s), .y(y2) );
  or_2_423 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_258 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_290 inv ( .a(s), .y(sa) );
  and_2_867 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_866 and2 ( .a(b), .b(s), .y(y2) );
  or_2_422 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_257 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_289 inv ( .a(s), .y(sa) );
  and_2_865 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_864 and2 ( .a(b), .b(s), .y(y2) );
  or_2_421 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_256 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_288 inv ( .a(s), .y(sa) );
  and_2_863 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_862 and2 ( .a(b), .b(s), .y(y2) );
  or_2_420 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_255 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_287 inv ( .a(s), .y(sa) );
  and_2_861 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_860 and2 ( .a(b), .b(s), .y(y2) );
  or_2_419 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_254 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_286 inv ( .a(s), .y(sa) );
  and_2_859 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_858 and2 ( .a(b), .b(s), .y(y2) );
  or_2_418 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_253 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_285 inv ( .a(s), .y(sa) );
  and_2_857 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_856 and2 ( .a(b), .b(s), .y(y2) );
  or_2_417 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_252 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_284 inv ( .a(s), .y(sa) );
  and_2_855 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_854 and2 ( .a(b), .b(s), .y(y2) );
  or_2_416 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_251 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_283 inv ( .a(s), .y(sa) );
  and_2_853 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_852 and2 ( .a(b), .b(s), .y(y2) );
  or_2_415 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_250 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_282 inv ( .a(s), .y(sa) );
  and_2_851 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_850 and2 ( .a(b), .b(s), .y(y2) );
  or_2_414 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_249 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_281 inv ( .a(s), .y(sa) );
  and_2_849 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_848 and2 ( .a(b), .b(s), .y(y2) );
  or_2_413 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_248 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_280 inv ( .a(s), .y(sa) );
  and_2_847 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_846 and2 ( .a(b), .b(s), .y(y2) );
  or_2_412 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_247 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_279 inv ( .a(s), .y(sa) );
  and_2_845 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_844 and2 ( .a(b), .b(s), .y(y2) );
  or_2_411 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_246 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_278 inv ( .a(s), .y(sa) );
  and_2_843 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_842 and2 ( .a(b), .b(s), .y(y2) );
  or_2_410 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_245 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_277 inv ( .a(s), .y(sa) );
  and_2_841 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_840 and2 ( .a(b), .b(s), .y(y2) );
  or_2_409 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_244 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_276 inv ( .a(s), .y(sa) );
  and_2_839 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_838 and2 ( .a(b), .b(s), .y(y2) );
  or_2_408 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_243 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_275 inv ( .a(s), .y(sa) );
  and_2_837 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_836 and2 ( .a(b), .b(s), .y(y2) );
  or_2_407 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_242 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_274 inv ( .a(s), .y(sa) );
  and_2_835 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_834 and2 ( .a(b), .b(s), .y(y2) );
  or_2_406 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_241 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_273 inv ( .a(s), .y(sa) );
  and_2_833 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_832 and2 ( .a(b), .b(s), .y(y2) );
  or_2_405 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_240 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_272 inv ( .a(s), .y(sa) );
  and_2_831 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_830 and2 ( .a(b), .b(s), .y(y2) );
  or_2_404 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_239 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_271 inv ( .a(s), .y(sa) );
  and_2_829 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_828 and2 ( .a(b), .b(s), .y(y2) );
  or_2_403 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_238 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_270 inv ( .a(s), .y(sa) );
  and_2_827 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_826 and2 ( .a(b), .b(s), .y(y2) );
  or_2_402 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_237 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_269 inv ( .a(s), .y(sa) );
  and_2_825 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_824 and2 ( .a(b), .b(s), .y(y2) );
  or_2_401 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_236 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_268 inv ( .a(s), .y(sa) );
  and_2_823 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_822 and2 ( .a(b), .b(s), .y(y2) );
  or_2_400 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_235 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_267 inv ( .a(s), .y(sa) );
  and_2_821 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_820 and2 ( .a(b), .b(s), .y(y2) );
  or_2_399 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_234 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_266 inv ( .a(s), .y(sa) );
  and_2_819 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_818 and2 ( .a(b), .b(s), .y(y2) );
  or_2_398 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_233 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_265 inv ( .a(s), .y(sa) );
  and_2_817 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_816 and2 ( .a(b), .b(s), .y(y2) );
  or_2_397 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_232 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_264 inv ( .a(s), .y(sa) );
  and_2_815 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_814 and2 ( .a(b), .b(s), .y(y2) );
  or_2_396 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_231 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_263 inv ( .a(s), .y(sa) );
  and_2_813 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_812 and2 ( .a(b), .b(s), .y(y2) );
  or_2_395 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_230 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_262 inv ( .a(s), .y(sa) );
  and_2_811 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_810 and2 ( .a(b), .b(s), .y(y2) );
  or_2_394 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_229 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_261 inv ( .a(s), .y(sa) );
  and_2_809 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_808 and2 ( .a(b), .b(s), .y(y2) );
  or_2_393 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_228 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_260 inv ( .a(s), .y(sa) );
  and_2_807 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_806 and2 ( .a(b), .b(s), .y(y2) );
  or_2_392 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_227 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_259 inv ( .a(s), .y(sa) );
  and_2_805 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_804 and2 ( .a(b), .b(s), .y(y2) );
  or_2_391 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_226 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_258 inv ( .a(s), .y(sa) );
  and_2_803 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_802 and2 ( .a(b), .b(s), .y(y2) );
  or_2_390 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_225 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_257 inv ( .a(s), .y(sa) );
  and_2_801 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_800 and2 ( .a(b), .b(s), .y(y2) );
  or_2_389 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_224 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_256 inv ( .a(s), .y(sa) );
  and_2_799 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_798 and2 ( .a(b), .b(s), .y(y2) );
  or_2_388 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_223 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_255 inv ( .a(s), .y(sa) );
  and_2_797 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_796 and2 ( .a(b), .b(s), .y(y2) );
  or_2_387 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_222 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_254 inv ( .a(s), .y(sa) );
  and_2_795 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_794 and2 ( .a(b), .b(s), .y(y2) );
  or_2_386 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_221 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_253 inv ( .a(s), .y(sa) );
  and_2_793 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_792 and2 ( .a(b), .b(s), .y(y2) );
  or_2_385 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_220 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_252 inv ( .a(s), .y(sa) );
  and_2_791 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_790 and2 ( .a(b), .b(s), .y(y2) );
  or_2_384 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_219 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_251 inv ( .a(s), .y(sa) );
  and_2_789 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_788 and2 ( .a(b), .b(s), .y(y2) );
  or_2_383 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_218 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_250 inv ( .a(s), .y(sa) );
  and_2_787 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_786 and2 ( .a(b), .b(s), .y(y2) );
  or_2_382 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_217 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_249 inv ( .a(s), .y(sa) );
  and_2_785 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_784 and2 ( .a(b), .b(s), .y(y2) );
  or_2_381 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_216 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_248 inv ( .a(s), .y(sa) );
  and_2_783 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_782 and2 ( .a(b), .b(s), .y(y2) );
  or_2_380 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_215 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_247 inv ( .a(s), .y(sa) );
  and_2_781 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_780 and2 ( .a(b), .b(s), .y(y2) );
  or_2_379 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_214 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_246 inv ( .a(s), .y(sa) );
  and_2_779 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_778 and2 ( .a(b), .b(s), .y(y2) );
  or_2_378 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_213 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_245 inv ( .a(s), .y(sa) );
  and_2_777 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_776 and2 ( .a(b), .b(s), .y(y2) );
  or_2_377 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_212 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_244 inv ( .a(s), .y(sa) );
  and_2_775 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_774 and2 ( .a(b), .b(s), .y(y2) );
  or_2_376 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_211 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_243 inv ( .a(s), .y(sa) );
  and_2_773 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_772 and2 ( .a(b), .b(s), .y(y2) );
  or_2_375 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_210 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_242 inv ( .a(s), .y(sa) );
  and_2_771 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_770 and2 ( .a(b), .b(s), .y(y2) );
  or_2_374 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_209 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_241 inv ( .a(s), .y(sa) );
  and_2_769 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_768 and2 ( .a(b), .b(s), .y(y2) );
  or_2_373 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_208 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_240 inv ( .a(s), .y(sa) );
  and_2_767 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_766 and2 ( .a(b), .b(s), .y(y2) );
  or_2_372 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_207 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_239 inv ( .a(s), .y(sa) );
  and_2_765 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_764 and2 ( .a(b), .b(s), .y(y2) );
  or_2_371 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_206 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_238 inv ( .a(s), .y(sa) );
  and_2_763 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_762 and2 ( .a(b), .b(s), .y(y2) );
  or_2_370 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_205 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_237 inv ( .a(s), .y(sa) );
  and_2_761 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_760 and2 ( .a(b), .b(s), .y(y2) );
  or_2_369 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_204 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_236 inv ( .a(s), .y(sa) );
  and_2_759 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_758 and2 ( .a(b), .b(s), .y(y2) );
  or_2_368 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_203 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_235 inv ( .a(s), .y(sa) );
  and_2_757 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_756 and2 ( .a(b), .b(s), .y(y2) );
  or_2_367 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_202 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_234 inv ( .a(s), .y(sa) );
  and_2_755 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_754 and2 ( .a(b), .b(s), .y(y2) );
  or_2_366 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_201 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_233 inv ( .a(s), .y(sa) );
  and_2_753 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_752 and2 ( .a(b), .b(s), .y(y2) );
  or_2_365 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_200 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_232 inv ( .a(s), .y(sa) );
  and_2_751 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_750 and2 ( .a(b), .b(s), .y(y2) );
  or_2_364 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_199 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_231 inv ( .a(s), .y(sa) );
  and_2_749 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_748 and2 ( .a(b), .b(s), .y(y2) );
  or_2_363 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_198 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_230 inv ( .a(s), .y(sa) );
  and_2_747 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_746 and2 ( .a(b), .b(s), .y(y2) );
  or_2_362 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_197 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_229 inv ( .a(s), .y(sa) );
  and_2_745 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_744 and2 ( .a(b), .b(s), .y(y2) );
  or_2_361 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_196 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_228 inv ( .a(s), .y(sa) );
  and_2_743 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_742 and2 ( .a(b), .b(s), .y(y2) );
  or_2_360 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_195 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_227 inv ( .a(s), .y(sa) );
  and_2_741 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_740 and2 ( .a(b), .b(s), .y(y2) );
  or_2_359 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_194 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_226 inv ( .a(s), .y(sa) );
  and_2_739 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_738 and2 ( .a(b), .b(s), .y(y2) );
  or_2_358 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_193 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_225 inv ( .a(s), .y(sa) );
  and_2_737 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_736 and2 ( .a(b), .b(s), .y(y2) );
  or_2_357 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_192 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_224 inv ( .a(s), .y(sa) );
  and_2_735 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_734 and2 ( .a(b), .b(s), .y(y2) );
  or_2_356 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_191 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_223 inv ( .a(s), .y(sa) );
  and_2_733 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_732 and2 ( .a(b), .b(s), .y(y2) );
  or_2_355 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_190 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_222 inv ( .a(s), .y(sa) );
  and_2_731 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_730 and2 ( .a(b), .b(s), .y(y2) );
  or_2_354 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_189 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_221 inv ( .a(s), .y(sa) );
  and_2_729 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_728 and2 ( .a(b), .b(s), .y(y2) );
  or_2_353 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_188 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_220 inv ( .a(s), .y(sa) );
  and_2_727 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_726 and2 ( .a(b), .b(s), .y(y2) );
  or_2_352 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_187 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_219 inv ( .a(s), .y(sa) );
  and_2_725 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_724 and2 ( .a(b), .b(s), .y(y2) );
  or_2_351 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_186 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_218 inv ( .a(s), .y(sa) );
  and_2_723 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_722 and2 ( .a(b), .b(s), .y(y2) );
  or_2_350 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_185 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_217 inv ( .a(s), .y(sa) );
  and_2_721 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_720 and2 ( .a(b), .b(s), .y(y2) );
  or_2_349 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_184 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_216 inv ( .a(s), .y(sa) );
  and_2_719 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_718 and2 ( .a(b), .b(s), .y(y2) );
  or_2_348 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_183 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_215 inv ( .a(s), .y(sa) );
  and_2_717 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_716 and2 ( .a(b), .b(s), .y(y2) );
  or_2_347 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_182 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_214 inv ( .a(s), .y(sa) );
  and_2_715 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_714 and2 ( .a(b), .b(s), .y(y2) );
  or_2_346 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_181 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_213 inv ( .a(s), .y(sa) );
  and_2_713 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_712 and2 ( .a(b), .b(s), .y(y2) );
  or_2_345 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_180 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_212 inv ( .a(s), .y(sa) );
  and_2_711 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_710 and2 ( .a(b), .b(s), .y(y2) );
  or_2_344 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_179 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_211 inv ( .a(s), .y(sa) );
  and_2_709 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_708 and2 ( .a(b), .b(s), .y(y2) );
  or_2_343 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_178 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_210 inv ( .a(s), .y(sa) );
  and_2_707 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_706 and2 ( .a(b), .b(s), .y(y2) );
  or_2_342 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_177 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_209 inv ( .a(s), .y(sa) );
  and_2_705 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_704 and2 ( .a(b), .b(s), .y(y2) );
  or_2_341 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_176 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_208 inv ( .a(s), .y(sa) );
  and_2_703 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_702 and2 ( .a(b), .b(s), .y(y2) );
  or_2_340 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_175 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_207 inv ( .a(s), .y(sa) );
  and_2_701 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_700 and2 ( .a(b), .b(s), .y(y2) );
  or_2_339 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_174 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_206 inv ( .a(s), .y(sa) );
  and_2_699 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_698 and2 ( .a(b), .b(s), .y(y2) );
  or_2_338 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_173 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_205 inv ( .a(s), .y(sa) );
  and_2_697 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_696 and2 ( .a(b), .b(s), .y(y2) );
  or_2_337 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_172 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_204 inv ( .a(s), .y(sa) );
  and_2_695 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_694 and2 ( .a(b), .b(s), .y(y2) );
  or_2_336 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_171 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_203 inv ( .a(s), .y(sa) );
  and_2_693 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_692 and2 ( .a(b), .b(s), .y(y2) );
  or_2_335 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_170 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_202 inv ( .a(s), .y(sa) );
  and_2_691 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_690 and2 ( .a(b), .b(s), .y(y2) );
  or_2_334 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_169 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_201 inv ( .a(s), .y(sa) );
  and_2_689 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_688 and2 ( .a(b), .b(s), .y(y2) );
  or_2_333 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_168 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_200 inv ( .a(s), .y(sa) );
  and_2_687 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_686 and2 ( .a(b), .b(s), .y(y2) );
  or_2_332 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_167 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_199 inv ( .a(s), .y(sa) );
  and_2_685 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_684 and2 ( .a(b), .b(s), .y(y2) );
  or_2_331 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_166 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_198 inv ( .a(s), .y(sa) );
  and_2_683 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_682 and2 ( .a(b), .b(s), .y(y2) );
  or_2_330 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_165 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_197 inv ( .a(s), .y(sa) );
  and_2_681 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_680 and2 ( .a(b), .b(s), .y(y2) );
  or_2_329 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_164 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_196 inv ( .a(s), .y(sa) );
  and_2_679 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_678 and2 ( .a(b), .b(s), .y(y2) );
  or_2_328 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_163 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_195 inv ( .a(s), .y(sa) );
  and_2_677 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_676 and2 ( .a(b), .b(s), .y(y2) );
  or_2_327 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_162 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_194 inv ( .a(s), .y(sa) );
  and_2_675 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_674 and2 ( .a(b), .b(s), .y(y2) );
  or_2_326 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_161 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_193 inv ( .a(s), .y(sa) );
  and_2_673 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_672 and2 ( .a(b), .b(s), .y(y2) );
  or_2_325 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_160 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_192 inv ( .a(s), .y(sa) );
  and_2_671 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_670 and2 ( .a(b), .b(s), .y(y2) );
  or_2_324 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_159 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_191 inv ( .a(s), .y(sa) );
  and_2_669 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_668 and2 ( .a(b), .b(s), .y(y2) );
  or_2_323 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_158 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_190 inv ( .a(s), .y(sa) );
  and_2_667 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_666 and2 ( .a(b), .b(s), .y(y2) );
  or_2_322 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_157 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_189 inv ( .a(s), .y(sa) );
  and_2_665 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_664 and2 ( .a(b), .b(s), .y(y2) );
  or_2_321 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_156 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_188 inv ( .a(s), .y(sa) );
  and_2_663 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_662 and2 ( .a(b), .b(s), .y(y2) );
  or_2_320 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_155 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_187 inv ( .a(s), .y(sa) );
  and_2_661 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_660 and2 ( .a(b), .b(s), .y(y2) );
  or_2_319 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_154 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_186 inv ( .a(s), .y(sa) );
  and_2_659 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_658 and2 ( .a(b), .b(s), .y(y2) );
  or_2_318 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_153 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_185 inv ( .a(s), .y(sa) );
  and_2_657 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_656 and2 ( .a(b), .b(s), .y(y2) );
  or_2_317 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_152 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_184 inv ( .a(s), .y(sa) );
  and_2_655 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_654 and2 ( .a(b), .b(s), .y(y2) );
  or_2_316 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_151 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_183 inv ( .a(s), .y(sa) );
  and_2_653 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_652 and2 ( .a(b), .b(s), .y(y2) );
  or_2_315 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_150 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_182 inv ( .a(s), .y(sa) );
  and_2_651 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_650 and2 ( .a(b), .b(s), .y(y2) );
  or_2_314 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_149 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_181 inv ( .a(s), .y(sa) );
  and_2_649 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_648 and2 ( .a(b), .b(s), .y(y2) );
  or_2_313 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_148 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_180 inv ( .a(s), .y(sa) );
  and_2_647 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_646 and2 ( .a(b), .b(s), .y(y2) );
  or_2_312 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_147 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_179 inv ( .a(s), .y(sa) );
  and_2_645 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_644 and2 ( .a(b), .b(s), .y(y2) );
  or_2_311 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_146 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_178 inv ( .a(s), .y(sa) );
  and_2_643 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_642 and2 ( .a(b), .b(s), .y(y2) );
  or_2_310 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_145 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_177 inv ( .a(s), .y(sa) );
  and_2_641 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_640 and2 ( .a(b), .b(s), .y(y2) );
  or_2_309 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_144 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_176 inv ( .a(s), .y(sa) );
  and_2_639 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_638 and2 ( .a(b), .b(s), .y(y2) );
  or_2_308 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_143 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_175 inv ( .a(s), .y(sa) );
  and_2_637 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_636 and2 ( .a(b), .b(s), .y(y2) );
  or_2_307 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_142 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_174 inv ( .a(s), .y(sa) );
  and_2_635 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_634 and2 ( .a(b), .b(s), .y(y2) );
  or_2_306 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_141 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_173 inv ( .a(s), .y(sa) );
  and_2_633 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_632 and2 ( .a(b), .b(s), .y(y2) );
  or_2_305 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_140 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_172 inv ( .a(s), .y(sa) );
  and_2_631 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_630 and2 ( .a(b), .b(s), .y(y2) );
  or_2_304 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_139 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_171 inv ( .a(s), .y(sa) );
  and_2_629 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_628 and2 ( .a(b), .b(s), .y(y2) );
  or_2_303 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_138 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_170 inv ( .a(s), .y(sa) );
  and_2_627 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_626 and2 ( .a(b), .b(s), .y(y2) );
  or_2_302 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_137 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_169 inv ( .a(s), .y(sa) );
  and_2_625 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_624 and2 ( .a(b), .b(s), .y(y2) );
  or_2_301 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_136 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_168 inv ( .a(s), .y(sa) );
  and_2_623 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_622 and2 ( .a(b), .b(s), .y(y2) );
  or_2_300 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_135 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_167 inv ( .a(s), .y(sa) );
  and_2_621 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_620 and2 ( .a(b), .b(s), .y(y2) );
  or_2_299 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_134 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_166 inv ( .a(s), .y(sa) );
  and_2_619 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_618 and2 ( .a(b), .b(s), .y(y2) );
  or_2_298 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_133 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_165 inv ( .a(s), .y(sa) );
  and_2_617 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_616 and2 ( .a(b), .b(s), .y(y2) );
  or_2_297 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_132 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_164 inv ( .a(s), .y(sa) );
  and_2_615 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_614 and2 ( .a(b), .b(s), .y(y2) );
  or_2_296 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_131 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_163 inv ( .a(s), .y(sa) );
  and_2_613 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_612 and2 ( .a(b), .b(s), .y(y2) );
  or_2_295 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_130 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_162 inv ( .a(s), .y(sa) );
  and_2_611 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_610 and2 ( .a(b), .b(s), .y(y2) );
  or_2_294 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_129 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_161 inv ( .a(s), .y(sa) );
  and_2_609 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_608 and2 ( .a(b), .b(s), .y(y2) );
  or_2_293 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_128 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_160 inv ( .a(s), .y(sa) );
  and_2_607 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_606 and2 ( .a(b), .b(s), .y(y2) );
  or_2_292 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_127 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_159 inv ( .a(s), .y(sa) );
  and_2_605 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_604 and2 ( .a(b), .b(s), .y(y2) );
  or_2_291 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_126 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_158 inv ( .a(s), .y(sa) );
  and_2_603 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_602 and2 ( .a(b), .b(s), .y(y2) );
  or_2_290 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_125 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_157 inv ( .a(s), .y(sa) );
  and_2_601 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_600 and2 ( .a(b), .b(s), .y(y2) );
  or_2_289 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_124 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_156 inv ( .a(s), .y(sa) );
  and_2_599 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_598 and2 ( .a(b), .b(s), .y(y2) );
  or_2_288 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_123 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_155 inv ( .a(s), .y(sa) );
  and_2_597 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_596 and2 ( .a(b), .b(s), .y(y2) );
  or_2_287 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_122 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_154 inv ( .a(s), .y(sa) );
  and_2_595 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_594 and2 ( .a(b), .b(s), .y(y2) );
  or_2_286 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_121 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_153 inv ( .a(s), .y(sa) );
  and_2_593 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_592 and2 ( .a(b), .b(s), .y(y2) );
  or_2_285 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_120 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_152 inv ( .a(s), .y(sa) );
  and_2_591 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_590 and2 ( .a(b), .b(s), .y(y2) );
  or_2_284 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_119 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_151 inv ( .a(s), .y(sa) );
  and_2_589 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_588 and2 ( .a(b), .b(s), .y(y2) );
  or_2_283 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_118 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_150 inv ( .a(s), .y(sa) );
  and_2_587 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_586 and2 ( .a(b), .b(s), .y(y2) );
  or_2_282 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_117 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_149 inv ( .a(s), .y(sa) );
  and_2_585 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_584 and2 ( .a(b), .b(s), .y(y2) );
  or_2_281 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_116 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_148 inv ( .a(s), .y(sa) );
  and_2_583 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_582 and2 ( .a(b), .b(s), .y(y2) );
  or_2_280 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_115 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_147 inv ( .a(s), .y(sa) );
  and_2_581 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_580 and2 ( .a(b), .b(s), .y(y2) );
  or_2_279 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_114 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_146 inv ( .a(s), .y(sa) );
  and_2_579 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_578 and2 ( .a(b), .b(s), .y(y2) );
  or_2_278 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_113 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_145 inv ( .a(s), .y(sa) );
  and_2_577 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_576 and2 ( .a(b), .b(s), .y(y2) );
  or_2_277 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_112 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_144 inv ( .a(s), .y(sa) );
  and_2_575 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_574 and2 ( .a(b), .b(s), .y(y2) );
  or_2_276 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_111 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_143 inv ( .a(s), .y(sa) );
  and_2_573 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_572 and2 ( .a(b), .b(s), .y(y2) );
  or_2_275 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_110 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_142 inv ( .a(s), .y(sa) );
  and_2_571 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_570 and2 ( .a(b), .b(s), .y(y2) );
  or_2_274 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_109 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_141 inv ( .a(s), .y(sa) );
  and_2_569 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_568 and2 ( .a(b), .b(s), .y(y2) );
  or_2_273 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_108 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_140 inv ( .a(s), .y(sa) );
  and_2_567 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_566 and2 ( .a(b), .b(s), .y(y2) );
  or_2_272 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_107 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_139 inv ( .a(s), .y(sa) );
  and_2_565 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_564 and2 ( .a(b), .b(s), .y(y2) );
  or_2_271 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_106 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_138 inv ( .a(s), .y(sa) );
  and_2_563 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_562 and2 ( .a(b), .b(s), .y(y2) );
  or_2_270 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_105 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_137 inv ( .a(s), .y(sa) );
  and_2_561 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_560 and2 ( .a(b), .b(s), .y(y2) );
  or_2_269 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_104 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_136 inv ( .a(s), .y(sa) );
  and_2_559 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_558 and2 ( .a(b), .b(s), .y(y2) );
  or_2_268 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_103 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_135 inv ( .a(s), .y(sa) );
  and_2_557 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_556 and2 ( .a(b), .b(s), .y(y2) );
  or_2_267 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_102 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_134 inv ( .a(s), .y(sa) );
  and_2_555 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_554 and2 ( .a(b), .b(s), .y(y2) );
  or_2_266 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_101 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_133 inv ( .a(s), .y(sa) );
  and_2_553 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_552 and2 ( .a(b), .b(s), .y(y2) );
  or_2_265 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_100 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_132 inv ( .a(s), .y(sa) );
  and_2_551 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_550 and2 ( .a(b), .b(s), .y(y2) );
  or_2_264 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_99 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_131 inv ( .a(s), .y(sa) );
  and_2_549 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_548 and2 ( .a(b), .b(s), .y(y2) );
  or_2_263 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_98 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_130 inv ( .a(s), .y(sa) );
  and_2_547 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_546 and2 ( .a(b), .b(s), .y(y2) );
  or_2_262 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_97 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_129 inv ( .a(s), .y(sa) );
  and_2_545 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_544 and2 ( .a(b), .b(s), .y(y2) );
  or_2_261 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_96 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_128 inv ( .a(s), .y(sa) );
  and_2_543 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_542 and2 ( .a(b), .b(s), .y(y2) );
  or_2_260 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_95 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_127 inv ( .a(s), .y(sa) );
  and_2_541 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_540 and2 ( .a(b), .b(s), .y(y2) );
  or_2_259 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_94 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_126 inv ( .a(s), .y(sa) );
  and_2_539 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_538 and2 ( .a(b), .b(s), .y(y2) );
  or_2_258 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_93 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_125 inv ( .a(s), .y(sa) );
  and_2_537 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_536 and2 ( .a(b), .b(s), .y(y2) );
  or_2_257 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_92 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_124 inv ( .a(s), .y(sa) );
  and_2_535 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_534 and2 ( .a(b), .b(s), .y(y2) );
  or_2_256 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_91 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_123 inv ( .a(s), .y(sa) );
  and_2_533 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_532 and2 ( .a(b), .b(s), .y(y2) );
  or_2_255 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_90 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_122 inv ( .a(s), .y(sa) );
  and_2_531 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_530 and2 ( .a(b), .b(s), .y(y2) );
  or_2_254 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_89 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_121 inv ( .a(s), .y(sa) );
  and_2_529 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_528 and2 ( .a(b), .b(s), .y(y2) );
  or_2_253 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_88 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_120 inv ( .a(s), .y(sa) );
  and_2_527 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_526 and2 ( .a(b), .b(s), .y(y2) );
  or_2_252 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_87 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_119 inv ( .a(s), .y(sa) );
  and_2_525 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_524 and2 ( .a(b), .b(s), .y(y2) );
  or_2_251 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_86 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_118 inv ( .a(s), .y(sa) );
  and_2_523 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_522 and2 ( .a(b), .b(s), .y(y2) );
  or_2_250 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_85 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_117 inv ( .a(s), .y(sa) );
  and_2_521 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_520 and2 ( .a(b), .b(s), .y(y2) );
  or_2_249 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_84 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_116 inv ( .a(s), .y(sa) );
  and_2_519 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_518 and2 ( .a(b), .b(s), .y(y2) );
  or_2_248 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_83 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_115 inv ( .a(s), .y(sa) );
  and_2_517 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_516 and2 ( .a(b), .b(s), .y(y2) );
  or_2_247 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_82 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_114 inv ( .a(s), .y(sa) );
  and_2_515 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_514 and2 ( .a(b), .b(s), .y(y2) );
  or_2_246 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_81 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_113 inv ( .a(s), .y(sa) );
  and_2_513 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_512 and2 ( .a(b), .b(s), .y(y2) );
  or_2_245 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_80 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_112 inv ( .a(s), .y(sa) );
  and_2_511 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_510 and2 ( .a(b), .b(s), .y(y2) );
  or_2_244 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_79 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_111 inv ( .a(s), .y(sa) );
  and_2_509 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_508 and2 ( .a(b), .b(s), .y(y2) );
  or_2_243 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_78 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_110 inv ( .a(s), .y(sa) );
  and_2_507 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_506 and2 ( .a(b), .b(s), .y(y2) );
  or_2_242 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_77 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_109 inv ( .a(s), .y(sa) );
  and_2_505 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_504 and2 ( .a(b), .b(s), .y(y2) );
  or_2_241 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_76 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_108 inv ( .a(s), .y(sa) );
  and_2_503 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_502 and2 ( .a(b), .b(s), .y(y2) );
  or_2_240 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_75 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_107 inv ( .a(s), .y(sa) );
  and_2_501 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_500 and2 ( .a(b), .b(s), .y(y2) );
  or_2_239 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_74 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_106 inv ( .a(s), .y(sa) );
  and_2_499 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_498 and2 ( .a(b), .b(s), .y(y2) );
  or_2_238 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_73 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_105 inv ( .a(s), .y(sa) );
  and_2_497 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_496 and2 ( .a(b), .b(s), .y(y2) );
  or_2_237 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_72 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_104 inv ( .a(s), .y(sa) );
  and_2_495 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_494 and2 ( .a(b), .b(s), .y(y2) );
  or_2_236 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_71 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_103 inv ( .a(s), .y(sa) );
  and_2_493 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_492 and2 ( .a(b), .b(s), .y(y2) );
  or_2_235 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_70 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_102 inv ( .a(s), .y(sa) );
  and_2_491 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_490 and2 ( .a(b), .b(s), .y(y2) );
  or_2_234 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_69 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_101 inv ( .a(s), .y(sa) );
  and_2_489 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_488 and2 ( .a(b), .b(s), .y(y2) );
  or_2_233 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_68 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_100 inv ( .a(s), .y(sa) );
  and_2_487 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_486 and2 ( .a(b), .b(s), .y(y2) );
  or_2_232 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_67 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_99 inv ( .a(s), .y(sa) );
  and_2_485 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_484 and2 ( .a(b), .b(s), .y(y2) );
  or_2_231 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_66 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_98 inv ( .a(s), .y(sa) );
  and_2_483 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_482 and2 ( .a(b), .b(s), .y(y2) );
  or_2_230 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_65 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_97 inv ( .a(s), .y(sa) );
  and_2_481 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_480 and2 ( .a(b), .b(s), .y(y2) );
  or_2_229 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_64 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_96 inv ( .a(s), .y(sa) );
  and_2_479 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_478 and2 ( .a(b), .b(s), .y(y2) );
  or_2_228 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_63 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_95 inv ( .a(s), .y(sa) );
  and_2_477 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_476 and2 ( .a(b), .b(s), .y(y2) );
  or_2_227 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_62 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_94 inv ( .a(s), .y(sa) );
  and_2_475 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_474 and2 ( .a(b), .b(s), .y(y2) );
  or_2_226 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_61 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_93 inv ( .a(s), .y(sa) );
  and_2_473 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_472 and2 ( .a(b), .b(s), .y(y2) );
  or_2_225 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_60 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_92 inv ( .a(s), .y(sa) );
  and_2_471 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_470 and2 ( .a(b), .b(s), .y(y2) );
  or_2_224 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_59 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_91 inv ( .a(s), .y(sa) );
  and_2_469 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_468 and2 ( .a(b), .b(s), .y(y2) );
  or_2_223 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_58 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_90 inv ( .a(s), .y(sa) );
  and_2_467 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_466 and2 ( .a(b), .b(s), .y(y2) );
  or_2_222 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_57 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_89 inv ( .a(s), .y(sa) );
  and_2_465 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_464 and2 ( .a(b), .b(s), .y(y2) );
  or_2_221 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_56 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_88 inv ( .a(s), .y(sa) );
  and_2_463 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_462 and2 ( .a(b), .b(s), .y(y2) );
  or_2_220 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_55 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_87 inv ( .a(s), .y(sa) );
  and_2_461 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_460 and2 ( .a(b), .b(s), .y(y2) );
  or_2_219 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_54 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_86 inv ( .a(s), .y(sa) );
  and_2_459 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_458 and2 ( .a(b), .b(s), .y(y2) );
  or_2_218 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_53 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_85 inv ( .a(s), .y(sa) );
  and_2_457 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_456 and2 ( .a(b), .b(s), .y(y2) );
  or_2_217 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_52 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_84 inv ( .a(s), .y(sa) );
  and_2_455 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_454 and2 ( .a(b), .b(s), .y(y2) );
  or_2_216 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_51 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_83 inv ( .a(s), .y(sa) );
  and_2_453 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_452 and2 ( .a(b), .b(s), .y(y2) );
  or_2_215 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_50 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_82 inv ( .a(s), .y(sa) );
  and_2_451 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_450 and2 ( .a(b), .b(s), .y(y2) );
  or_2_214 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_49 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_81 inv ( .a(s), .y(sa) );
  and_2_449 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_448 and2 ( .a(b), .b(s), .y(y2) );
  or_2_213 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_48 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_80 inv ( .a(s), .y(sa) );
  and_2_447 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_446 and2 ( .a(b), .b(s), .y(y2) );
  or_2_212 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_47 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_79 inv ( .a(s), .y(sa) );
  and_2_445 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_444 and2 ( .a(b), .b(s), .y(y2) );
  or_2_211 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_46 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_78 inv ( .a(s), .y(sa) );
  and_2_443 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_442 and2 ( .a(b), .b(s), .y(y2) );
  or_2_210 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_45 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_77 inv ( .a(s), .y(sa) );
  and_2_441 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_440 and2 ( .a(b), .b(s), .y(y2) );
  or_2_209 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_44 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_76 inv ( .a(s), .y(sa) );
  and_2_439 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_438 and2 ( .a(b), .b(s), .y(y2) );
  or_2_208 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_43 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_75 inv ( .a(s), .y(sa) );
  and_2_437 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_436 and2 ( .a(b), .b(s), .y(y2) );
  or_2_207 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_42 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_74 inv ( .a(s), .y(sa) );
  and_2_435 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_434 and2 ( .a(b), .b(s), .y(y2) );
  or_2_206 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_41 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_73 inv ( .a(s), .y(sa) );
  and_2_433 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_432 and2 ( .a(b), .b(s), .y(y2) );
  or_2_205 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_40 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_72 inv ( .a(s), .y(sa) );
  and_2_431 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_430 and2 ( .a(b), .b(s), .y(y2) );
  or_2_204 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_39 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_71 inv ( .a(s), .y(sa) );
  and_2_429 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_428 and2 ( .a(b), .b(s), .y(y2) );
  or_2_203 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_38 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_70 inv ( .a(s), .y(sa) );
  and_2_427 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_426 and2 ( .a(b), .b(s), .y(y2) );
  or_2_202 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_37 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_69 inv ( .a(s), .y(sa) );
  and_2_425 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_424 and2 ( .a(b), .b(s), .y(y2) );
  or_2_201 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_36 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_68 inv ( .a(s), .y(sa) );
  and_2_423 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_422 and2 ( .a(b), .b(s), .y(y2) );
  or_2_200 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_35 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_67 inv ( .a(s), .y(sa) );
  and_2_421 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_420 and2 ( .a(b), .b(s), .y(y2) );
  or_2_199 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_34 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_66 inv ( .a(s), .y(sa) );
  and_2_419 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_418 and2 ( .a(b), .b(s), .y(y2) );
  or_2_198 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_33 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;
  tri   y;

  not_1_65 inv ( .a(s), .y(sa) );
  and_2_417 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_416 and2 ( .a(b), .b(s), .y(y2) );
  or_2_197 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_32 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_32 inv ( .a(s), .y(sa) );
  and_2_176 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_175 and2 ( .a(b), .b(s), .y(y2) );
  or_2_88 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_31 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_31 inv ( .a(s), .y(sa) );
  and_2_174 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_173 and2 ( .a(b), .b(s), .y(y2) );
  or_2_87 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_30 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_30 inv ( .a(s), .y(sa) );
  and_2_172 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_171 and2 ( .a(b), .b(s), .y(y2) );
  or_2_86 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_29 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_29 inv ( .a(s), .y(sa) );
  and_2_170 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_169 and2 ( .a(b), .b(s), .y(y2) );
  or_2_85 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_28 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_28 inv ( .a(s), .y(sa) );
  and_2_152 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_151 and2 ( .a(b), .b(s), .y(y2) );
  or_2_76 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_27 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_27 inv ( .a(s), .y(sa) );
  and_2_150 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_149 and2 ( .a(b), .b(s), .y(y2) );
  or_2_75 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_26 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_26 inv ( .a(s), .y(sa) );
  and_2_148 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_147 and2 ( .a(b), .b(s), .y(y2) );
  or_2_74 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_25 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_25 inv ( .a(s), .y(sa) );
  and_2_146 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_145 and2 ( .a(b), .b(s), .y(y2) );
  or_2_73 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_24 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_24 inv ( .a(s), .y(sa) );
  and_2_128 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_127 and2 ( .a(b), .b(s), .y(y2) );
  or_2_64 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_23 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_23 inv ( .a(s), .y(sa) );
  and_2_126 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_125 and2 ( .a(b), .b(s), .y(y2) );
  or_2_63 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_22 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_22 inv ( .a(s), .y(sa) );
  and_2_124 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_123 and2 ( .a(b), .b(s), .y(y2) );
  or_2_62 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_21 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_21 inv ( .a(s), .y(sa) );
  and_2_122 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_121 and2 ( .a(b), .b(s), .y(y2) );
  or_2_61 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_20 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_20 inv ( .a(s), .y(sa) );
  and_2_104 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_103 and2 ( .a(b), .b(s), .y(y2) );
  or_2_52 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_19 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_19 inv ( .a(s), .y(sa) );
  and_2_102 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_101 and2 ( .a(b), .b(s), .y(y2) );
  or_2_51 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_18 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_18 inv ( .a(s), .y(sa) );
  and_2_100 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_99 and2 ( .a(b), .b(s), .y(y2) );
  or_2_50 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_17 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_17 inv ( .a(s), .y(sa) );
  and_2_98 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_97 and2 ( .a(b), .b(s), .y(y2) );
  or_2_49 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_16 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_16 inv ( .a(s), .y(sa) );
  and_2_80 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_79 and2 ( .a(b), .b(s), .y(y2) );
  or_2_40 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_15 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_15 inv ( .a(s), .y(sa) );
  and_2_78 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_77 and2 ( .a(b), .b(s), .y(y2) );
  or_2_39 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_14 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_14 inv ( .a(s), .y(sa) );
  and_2_76 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_75 and2 ( .a(b), .b(s), .y(y2) );
  or_2_38 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_13 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_13 inv ( .a(s), .y(sa) );
  and_2_74 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_73 and2 ( .a(b), .b(s), .y(y2) );
  or_2_37 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_12 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_12 inv ( .a(s), .y(sa) );
  and_2_56 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_55 and2 ( .a(b), .b(s), .y(y2) );
  or_2_28 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_11 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_11 inv ( .a(s), .y(sa) );
  and_2_54 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_53 and2 ( .a(b), .b(s), .y(y2) );
  or_2_27 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_10 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_10 inv ( .a(s), .y(sa) );
  and_2_52 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_51 and2 ( .a(b), .b(s), .y(y2) );
  or_2_26 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_9 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_9 inv ( .a(s), .y(sa) );
  and_2_50 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_49 and2 ( .a(b), .b(s), .y(y2) );
  or_2_25 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_8 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_8 inv ( .a(s), .y(sa) );
  and_2_32 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_31 and2 ( .a(b), .b(s), .y(y2) );
  or_2_16 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_7 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_7 inv ( .a(s), .y(sa) );
  and_2_30 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_29 and2 ( .a(b), .b(s), .y(y2) );
  or_2_15 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_6 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_6 inv ( .a(s), .y(sa) );
  and_2_28 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_27 and2 ( .a(b), .b(s), .y(y2) );
  or_2_14 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_5 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_5 inv ( .a(s), .y(sa) );
  and_2_26 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_25 and2 ( .a(b), .b(s), .y(y2) );
  or_2_13 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_4 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_4 inv ( .a(s), .y(sa) );
  and_2_8 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_7 and2 ( .a(b), .b(s), .y(y2) );
  or_2_4 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_3 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_3 inv ( .a(s), .y(sa) );
  and_2_6 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_5 and2 ( .a(b), .b(s), .y(y2) );
  or_2_3 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_2 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_2 inv ( .a(s), .y(sa) );
  and_2_4 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_3 and2 ( .a(b), .b(s), .y(y2) );
  or_2_2 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module mux21_1 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_1 inv ( .a(s), .y(sa) );
  and_2_2 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1 and2 ( .a(b), .b(s), .y(y2) );
  or_2_1 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module xnor_2_31 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_30 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_29 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_28 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_27 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_26 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_25 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_24 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_23 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_22 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_21 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_20 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_19 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_18 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_17 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_16 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_15 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_14 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_13 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_12 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_11 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_10 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_9 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_8 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_7 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_6 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_5 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_4 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_3 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_2 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module xnor_2_1 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module ffd_async_288 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_287 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_286 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_290 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;
  wire   n1;

  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q), .QN(n1) );
endmodule


module ffd_async_273 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;
  wire   n1;

  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q), .QN(n1) );
endmodule


module ffd_async_305 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_304 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_303 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_302 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_301 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_300 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_299 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_298 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_297 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_296 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_295 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_294 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_293 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_292 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_285 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_284 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_283 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_282 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_281 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_280 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_279 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_278 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_277 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_276 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_275 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_274 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_272 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_271 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_270 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_269 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_268 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_267 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_266 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_265 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_264 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_263 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_262 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_261 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_260 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_259 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_258 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_257 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_256 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_255 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_254 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_253 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_252 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_251 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_250 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_249 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_248 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_247 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_246 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_245 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_244 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_243 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_242 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_241 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_240 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_239 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_238 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_237 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_236 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_235 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_234 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_233 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_232 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_231 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_230 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_229 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_228 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_227 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_226 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_225 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_224 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_223 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_222 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_221 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_220 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_219 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_218 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_217 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_216 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_215 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_214 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_213 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_212 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_211 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_210 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_209 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_208 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_207 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_206 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_205 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_204 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_203 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_202 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_201 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_200 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_199 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_198 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_197 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_196 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_195 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_194 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_193 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_192 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_191 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_190 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_189 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_188 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_187 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_186 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_185 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_184 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_183 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_182 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_181 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_180 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_179 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_178 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_177 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_176 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_175 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_174 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_173 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_172 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_171 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_170 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_169 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_168 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_167 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_166 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_165 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_164 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_163 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_162 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_161 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_160 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_159 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_158 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_157 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_156 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_155 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_154 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_153 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_152 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_151 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_150 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_149 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_148 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_147 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_146 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_145 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_144 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_143 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_142 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_141 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_140 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_139 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_138 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_137 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_136 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_135 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_134 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_133 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_132 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_131 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_130 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_129 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_128 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_127 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_126 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_125 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_124 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_123 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_122 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_121 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_120 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_119 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_118 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_117 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_116 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_115 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_114 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_113 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_112 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_111 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_110 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_109 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_108 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_107 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_106 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_105 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_104 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_103 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_102 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_101 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_100 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_99 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_98 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_97 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_96 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_95 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_94 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_93 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_92 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_91 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_90 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_89 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_88 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_87 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_86 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_85 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_84 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_83 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_82 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_81 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_80 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_79 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_78 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_77 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_76 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_75 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_74 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_73 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_72 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_71 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_70 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_69 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_68 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_67 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_66 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_65 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_64 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_63 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_62 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_61 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_60 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_59 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_58 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_57 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_56 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_55 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_54 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_53 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_52 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_51 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_50 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_49 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_48 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_47 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_46 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_45 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_44 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_43 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_42 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_41 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_40 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_39 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_38 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_37 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_36 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_35 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_34 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_33 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_32 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_31 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_30 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_29 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_28 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_27 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_26 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_25 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_24 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_23 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_22 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_21 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_20 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_19 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_18 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_17 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_16 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_15 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_14 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_13 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_12 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_11 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_10 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_9 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_8 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_7 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_6 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_5 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_4 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_3 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_2 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_1 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module mux21_generic_n32_3 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n1, n2, n3;

  mux21_448 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(n1), .y(y[0]) );
  mux21_447 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(n1), .y(y[1]) );
  mux21_446 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(n1), .y(y[2]) );
  mux21_445 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(n1), .y(y[3]) );
  mux21_444 mux21_i_4 ( .a(a[4]), .b(b[4]), .s(n1), .y(y[4]) );
  mux21_443 mux21_i_5 ( .a(a[5]), .b(b[5]), .s(n1), .y(y[5]) );
  mux21_442 mux21_i_6 ( .a(a[6]), .b(b[6]), .s(n1), .y(y[6]) );
  mux21_441 mux21_i_7 ( .a(a[7]), .b(b[7]), .s(n1), .y(y[7]) );
  mux21_440 mux21_i_8 ( .a(a[8]), .b(b[8]), .s(n1), .y(y[8]) );
  mux21_439 mux21_i_9 ( .a(a[9]), .b(b[9]), .s(n1), .y(y[9]) );
  mux21_438 mux21_i_10 ( .a(a[10]), .b(b[10]), .s(n1), .y(y[10]) );
  mux21_437 mux21_i_11 ( .a(a[11]), .b(b[11]), .s(n1), .y(y[11]) );
  mux21_436 mux21_i_12 ( .a(a[12]), .b(b[12]), .s(n2), .y(y[12]) );
  mux21_435 mux21_i_13 ( .a(a[13]), .b(b[13]), .s(n2), .y(y[13]) );
  mux21_434 mux21_i_14 ( .a(a[14]), .b(b[14]), .s(n2), .y(y[14]) );
  mux21_433 mux21_i_15 ( .a(a[15]), .b(b[15]), .s(n2), .y(y[15]) );
  mux21_432 mux21_i_16 ( .a(a[16]), .b(b[16]), .s(n2), .y(y[16]) );
  mux21_431 mux21_i_17 ( .a(a[17]), .b(b[17]), .s(n2), .y(y[17]) );
  mux21_430 mux21_i_18 ( .a(a[18]), .b(b[18]), .s(n2), .y(y[18]) );
  mux21_429 mux21_i_19 ( .a(a[19]), .b(b[19]), .s(n2), .y(y[19]) );
  mux21_428 mux21_i_20 ( .a(a[20]), .b(b[20]), .s(n2), .y(y[20]) );
  mux21_427 mux21_i_21 ( .a(a[21]), .b(b[21]), .s(n2), .y(y[21]) );
  mux21_426 mux21_i_22 ( .a(a[22]), .b(b[22]), .s(n2), .y(y[22]) );
  mux21_425 mux21_i_23 ( .a(a[23]), .b(b[23]), .s(n2), .y(y[23]) );
  mux21_424 mux21_i_24 ( .a(a[24]), .b(b[24]), .s(n3), .y(y[24]) );
  mux21_423 mux21_i_25 ( .a(a[25]), .b(b[25]), .s(n3), .y(y[25]) );
  mux21_422 mux21_i_26 ( .a(a[26]), .b(b[26]), .s(n3), .y(y[26]) );
  mux21_421 mux21_i_27 ( .a(a[27]), .b(b[27]), .s(n3), .y(y[27]) );
  mux21_420 mux21_i_28 ( .a(a[28]), .b(b[28]), .s(n3), .y(y[28]) );
  mux21_419 mux21_i_29 ( .a(a[29]), .b(b[29]), .s(n3), .y(y[29]) );
  mux21_418 mux21_i_30 ( .a(a[30]), .b(b[30]), .s(n3), .y(y[30]) );
  mux21_417 mux21_i_31 ( .a(a[31]), .b(b[31]), .s(n3), .y(y[31]) );
  BUF_X1 U1 ( .A(sel), .Z(n1) );
  BUF_X1 U2 ( .A(sel), .Z(n2) );
  BUF_X1 U3 ( .A(sel), .Z(n3) );
endmodule


module mux21_generic_n32_2 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n1, n2, n3;

  mux21_416 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(n1), .y(y[0]) );
  mux21_415 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(n1), .y(y[1]) );
  mux21_414 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(n1), .y(y[2]) );
  mux21_413 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(n1), .y(y[3]) );
  mux21_412 mux21_i_4 ( .a(a[4]), .b(b[4]), .s(n1), .y(y[4]) );
  mux21_411 mux21_i_5 ( .a(a[5]), .b(b[5]), .s(n1), .y(y[5]) );
  mux21_410 mux21_i_6 ( .a(a[6]), .b(b[6]), .s(n1), .y(y[6]) );
  mux21_409 mux21_i_7 ( .a(a[7]), .b(b[7]), .s(n1), .y(y[7]) );
  mux21_408 mux21_i_8 ( .a(a[8]), .b(b[8]), .s(n1), .y(y[8]) );
  mux21_407 mux21_i_9 ( .a(a[9]), .b(b[9]), .s(n1), .y(y[9]) );
  mux21_406 mux21_i_10 ( .a(a[10]), .b(b[10]), .s(n1), .y(y[10]) );
  mux21_405 mux21_i_11 ( .a(a[11]), .b(b[11]), .s(n1), .y(y[11]) );
  mux21_404 mux21_i_12 ( .a(a[12]), .b(b[12]), .s(n2), .y(y[12]) );
  mux21_403 mux21_i_13 ( .a(a[13]), .b(b[13]), .s(n2), .y(y[13]) );
  mux21_402 mux21_i_14 ( .a(a[14]), .b(b[14]), .s(n2), .y(y[14]) );
  mux21_401 mux21_i_15 ( .a(a[15]), .b(b[15]), .s(n2), .y(y[15]) );
  mux21_400 mux21_i_16 ( .a(a[16]), .b(b[16]), .s(n2), .y(y[16]) );
  mux21_399 mux21_i_17 ( .a(a[17]), .b(b[17]), .s(n2), .y(y[17]) );
  mux21_398 mux21_i_18 ( .a(a[18]), .b(b[18]), .s(n2), .y(y[18]) );
  mux21_397 mux21_i_19 ( .a(a[19]), .b(b[19]), .s(n2), .y(y[19]) );
  mux21_396 mux21_i_20 ( .a(a[20]), .b(b[20]), .s(n2), .y(y[20]) );
  mux21_395 mux21_i_21 ( .a(a[21]), .b(b[21]), .s(n2), .y(y[21]) );
  mux21_394 mux21_i_22 ( .a(a[22]), .b(b[22]), .s(n2), .y(y[22]) );
  mux21_393 mux21_i_23 ( .a(a[23]), .b(b[23]), .s(n2), .y(y[23]) );
  mux21_392 mux21_i_24 ( .a(a[24]), .b(b[24]), .s(n3), .y(y[24]) );
  mux21_391 mux21_i_25 ( .a(a[25]), .b(b[25]), .s(n3), .y(y[25]) );
  mux21_390 mux21_i_26 ( .a(a[26]), .b(b[26]), .s(n3), .y(y[26]) );
  mux21_389 mux21_i_27 ( .a(a[27]), .b(b[27]), .s(n3), .y(y[27]) );
  mux21_388 mux21_i_28 ( .a(a[28]), .b(b[28]), .s(n3), .y(y[28]) );
  mux21_387 mux21_i_29 ( .a(a[29]), .b(b[29]), .s(n3), .y(y[29]) );
  mux21_386 mux21_i_30 ( .a(a[30]), .b(b[30]), .s(n3), .y(y[30]) );
  mux21_385 mux21_i_31 ( .a(a[31]), .b(b[31]), .s(n3), .y(y[31]) );
  BUF_X1 U1 ( .A(sel), .Z(n2) );
  BUF_X1 U2 ( .A(sel), .Z(n1) );
  BUF_X1 U3 ( .A(sel), .Z(n3) );
endmodule


module mux21_generic_n32_1 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n1, n2, n3;

  mux21_384 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(n1), .y(y[0]) );
  mux21_383 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(n1), .y(y[1]) );
  mux21_382 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(n1), .y(y[2]) );
  mux21_381 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(n1), .y(y[3]) );
  mux21_380 mux21_i_4 ( .a(a[4]), .b(b[4]), .s(n1), .y(y[4]) );
  mux21_379 mux21_i_5 ( .a(a[5]), .b(b[5]), .s(n1), .y(y[5]) );
  mux21_378 mux21_i_6 ( .a(a[6]), .b(b[6]), .s(n1), .y(y[6]) );
  mux21_377 mux21_i_7 ( .a(a[7]), .b(b[7]), .s(n1), .y(y[7]) );
  mux21_376 mux21_i_8 ( .a(a[8]), .b(b[8]), .s(n1), .y(y[8]) );
  mux21_375 mux21_i_9 ( .a(a[9]), .b(b[9]), .s(n1), .y(y[9]) );
  mux21_374 mux21_i_10 ( .a(a[10]), .b(b[10]), .s(n1), .y(y[10]) );
  mux21_373 mux21_i_11 ( .a(a[11]), .b(b[11]), .s(n1), .y(y[11]) );
  mux21_372 mux21_i_12 ( .a(a[12]), .b(b[12]), .s(n2), .y(y[12]) );
  mux21_371 mux21_i_13 ( .a(a[13]), .b(b[13]), .s(n2), .y(y[13]) );
  mux21_370 mux21_i_14 ( .a(a[14]), .b(b[14]), .s(n2), .y(y[14]) );
  mux21_369 mux21_i_15 ( .a(a[15]), .b(b[15]), .s(n2), .y(y[15]) );
  mux21_368 mux21_i_16 ( .a(a[16]), .b(b[16]), .s(n2), .y(y[16]) );
  mux21_367 mux21_i_17 ( .a(a[17]), .b(b[17]), .s(n2), .y(y[17]) );
  mux21_366 mux21_i_18 ( .a(a[18]), .b(b[18]), .s(n2), .y(y[18]) );
  mux21_365 mux21_i_19 ( .a(a[19]), .b(b[19]), .s(n2), .y(y[19]) );
  mux21_364 mux21_i_20 ( .a(a[20]), .b(b[20]), .s(n2), .y(y[20]) );
  mux21_363 mux21_i_21 ( .a(a[21]), .b(b[21]), .s(n2), .y(y[21]) );
  mux21_362 mux21_i_22 ( .a(a[22]), .b(b[22]), .s(n2), .y(y[22]) );
  mux21_361 mux21_i_23 ( .a(a[23]), .b(b[23]), .s(n2), .y(y[23]) );
  mux21_360 mux21_i_24 ( .a(a[24]), .b(b[24]), .s(n3), .y(y[24]) );
  mux21_359 mux21_i_25 ( .a(a[25]), .b(b[25]), .s(n3), .y(y[25]) );
  mux21_358 mux21_i_26 ( .a(a[26]), .b(b[26]), .s(n3), .y(y[26]) );
  mux21_357 mux21_i_27 ( .a(a[27]), .b(b[27]), .s(n3), .y(y[27]) );
  mux21_356 mux21_i_28 ( .a(a[28]), .b(b[28]), .s(n3), .y(y[28]) );
  mux21_355 mux21_i_29 ( .a(a[29]), .b(b[29]), .s(n3), .y(y[29]) );
  mux21_354 mux21_i_30 ( .a(a[30]), .b(b[30]), .s(n3), .y(y[30]) );
  mux21_353 mux21_i_31 ( .a(a[31]), .b(b[31]), .s(n3), .y(y[31]) );
  BUF_X1 U1 ( .A(sel), .Z(n1) );
  BUF_X1 U2 ( .A(sel), .Z(n2) );
  BUF_X1 U3 ( .A(sel), .Z(n3) );
endmodule


module and_2_1374 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1373 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1372 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1371 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1370 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1369 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1368 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1367 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1366 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1365 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1364 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1363 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1362 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1361 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1360 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1359 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1358 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1357 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1356 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1355 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1354 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1353 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1352 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1351 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1350 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1349 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1348 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1347 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1346 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1345 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1344 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1343 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1342 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1341 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1340 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1339 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1338 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1337 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1336 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1335 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1334 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1333 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1332 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1331 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1330 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1329 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1328 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1327 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1326 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1325 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1324 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1323 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1322 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1321 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1320 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1319 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1318 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1317 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1316 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1315 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1314 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1313 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1312 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1311 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1310 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1309 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1308 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1307 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1306 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1305 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1304 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1303 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1302 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1301 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1300 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1299 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1298 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1297 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1296 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1295 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1294 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1293 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1292 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1291 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1290 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1289 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1288 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1287 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1286 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1285 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1284 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1283 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1282 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1281 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1280 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1279 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1278 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1277 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1276 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1275 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1274 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1273 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1272 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1271 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1270 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1269 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1268 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1267 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1266 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1265 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1264 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1263 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1262 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1261 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1260 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1259 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1258 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1257 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1256 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1255 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1254 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1253 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1252 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1251 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1250 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1249 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1248 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1247 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1246 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1245 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1244 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1243 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1242 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1241 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1240 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1239 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1238 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1237 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1236 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1235 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1234 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1233 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1232 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1231 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1230 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1229 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1228 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1227 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1226 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1225 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1224 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1223 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1222 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1221 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1220 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1219 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1218 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1217 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1216 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1215 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1214 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1213 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1212 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1211 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1210 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1209 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1208 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1207 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1206 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1205 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1204 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1203 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1202 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1201 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1200 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1199 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1198 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1197 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1196 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1195 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1194 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1193 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1192 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1191 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1190 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1189 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1188 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1187 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1186 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1185 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1184 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1183 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1182 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1181 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1180 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1179 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1178 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1177 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1176 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1175 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1174 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1173 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1172 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1171 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1170 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1169 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1168 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1167 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1166 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1165 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1164 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1163 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1162 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1161 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1160 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1159 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1158 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1157 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1156 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1155 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1154 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1153 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1152 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1151 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1150 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1149 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1148 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1147 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1146 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1145 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1144 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1143 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1142 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1141 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1140 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1139 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1138 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1137 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1136 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1135 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1134 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1133 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1132 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1131 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1130 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1129 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1128 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1127 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1126 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1125 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1124 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1123 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1122 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1121 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1120 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1119 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1118 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1117 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1116 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1115 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1114 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1113 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1112 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1111 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1110 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1109 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1108 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1107 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1106 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1105 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1104 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1103 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1102 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1101 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1100 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1099 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1098 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1097 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1096 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1095 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1094 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1093 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1092 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1091 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1090 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1089 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1088 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1087 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1086 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1085 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1084 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1083 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1082 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1081 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1080 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1079 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1078 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1077 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1076 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1075 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1074 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1073 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1072 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1071 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1070 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1069 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1068 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1067 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1066 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1065 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1064 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1063 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1062 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1061 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1060 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1059 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1058 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1057 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1056 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1055 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1054 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1053 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1052 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1051 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1050 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1049 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1048 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1047 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1046 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1045 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1044 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1043 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1042 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1041 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1040 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1039 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1038 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1037 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1036 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1035 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1034 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1033 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1032 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1031 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1030 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1029 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1028 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1027 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1026 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1025 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1024 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1023 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1022 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1021 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1020 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1019 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1018 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1017 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1016 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1015 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1014 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1013 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1012 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1011 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1010 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1009 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1008 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1007 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1006 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1005 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1004 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1003 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1002 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1001 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1000 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_999 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_998 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_997 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_996 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_995 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_994 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_993 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_992 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_991 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_990 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_989 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_988 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_987 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_986 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_985 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_984 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_983 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_982 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_981 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_980 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_979 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_978 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_977 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_976 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_975 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_974 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_973 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_972 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_971 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_970 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_969 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_968 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_967 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_966 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_965 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_964 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_963 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_962 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_961 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_960 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_959 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_958 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_957 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_956 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_955 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_954 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_953 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_952 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_951 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_950 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_949 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_948 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_947 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_946 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_945 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_944 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_943 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_942 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_941 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_940 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_939 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_938 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_937 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_936 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_935 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_934 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_933 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_932 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_931 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_930 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_929 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_928 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_927 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_926 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_925 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_924 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_923 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_922 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_921 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_920 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_919 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_918 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_917 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_916 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_915 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_914 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_913 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_912 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_911 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_910 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_909 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_908 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_907 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_906 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_905 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_904 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_903 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_902 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_901 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_900 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_899 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_898 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_897 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_896 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_895 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_894 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_893 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_892 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_891 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_890 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_889 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_888 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_887 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_886 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_885 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_884 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_883 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_882 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_881 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_880 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_879 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_878 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_877 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_876 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_875 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_874 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_873 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_872 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_871 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_870 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_869 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_868 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_867 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_866 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_865 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_864 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_863 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_862 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_861 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_860 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_859 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_858 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_857 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_856 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_855 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_854 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_853 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_852 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_851 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_850 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_849 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_848 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_847 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_846 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_845 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_844 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_843 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_842 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_841 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_840 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_839 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_838 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_837 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_836 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_835 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_834 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_833 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_832 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_831 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_830 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_829 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_828 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_827 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_826 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_825 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_824 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_823 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_822 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_821 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_820 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_819 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_818 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_817 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_816 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_815 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_814 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_813 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_812 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_811 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_810 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_809 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_808 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_807 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_806 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_805 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_804 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_803 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_802 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_801 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_800 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_799 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_798 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_797 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_796 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_795 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_794 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_793 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_792 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_791 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_790 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_789 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_788 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_787 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_786 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_785 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_784 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_783 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_782 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_781 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_780 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_779 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_778 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_777 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_776 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_775 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_774 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_773 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_772 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_771 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_770 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_769 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_768 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_767 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_766 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_765 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_764 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_763 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_762 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_761 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_760 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_759 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_758 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_757 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_756 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_755 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_754 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_753 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_752 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_751 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_750 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_749 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_748 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_747 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_746 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_745 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_744 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_743 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_742 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_741 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_740 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_739 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_738 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_737 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_736 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_735 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_734 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_733 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_732 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_731 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_730 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_729 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_728 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_727 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_726 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_725 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_724 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_723 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_722 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_721 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_720 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_719 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_718 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_717 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_716 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_715 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_714 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_713 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_712 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_711 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_710 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_709 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_708 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_707 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_706 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_705 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_704 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_703 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_702 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_701 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_700 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_699 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_698 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_697 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_696 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_695 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_694 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_693 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_692 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_691 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_690 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_689 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_688 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_687 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_686 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_685 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_684 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_683 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_682 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_681 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_680 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_679 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_678 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_677 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_676 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_675 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_674 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_673 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_672 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_671 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_670 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_669 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_668 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_667 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_666 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_665 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_664 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_663 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_662 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_661 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_660 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_659 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_658 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_657 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_656 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_655 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_654 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_653 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_652 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_651 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_650 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_649 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_648 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_647 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_646 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_645 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_644 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_643 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_642 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_641 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_640 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_639 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_638 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_637 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_636 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_635 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_634 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_633 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_632 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_631 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_630 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_629 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_628 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_627 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_626 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_625 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_624 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_623 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_622 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_621 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_620 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_619 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_618 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_617 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_616 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_615 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_614 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_613 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_612 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_611 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_610 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_609 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_608 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_607 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_606 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_605 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_604 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_603 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_602 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_601 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_600 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_599 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_598 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_597 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_596 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_595 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_594 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_593 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_592 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_591 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_590 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_589 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_588 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_587 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_586 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_585 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_584 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_583 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_582 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_581 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_580 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_579 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_578 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_577 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_576 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_575 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_574 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_573 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_572 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_571 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_570 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_569 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_568 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_567 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_566 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_565 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_564 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_563 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_562 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_561 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_560 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_559 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_558 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_557 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_556 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_555 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_554 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_553 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_552 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_551 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_550 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_549 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_548 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_547 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_546 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_545 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_544 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_543 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_542 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_541 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_540 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_539 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_538 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_537 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_536 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_535 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_534 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_533 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_532 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_531 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_530 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_529 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_528 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_527 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_526 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_525 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_524 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_523 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_522 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_521 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_520 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_519 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_518 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_517 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_516 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_515 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_514 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_513 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_512 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_511 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_510 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_509 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_508 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_507 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_506 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_505 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_504 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_503 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_502 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_501 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_500 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_499 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_498 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_497 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_496 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_495 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_494 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_493 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_492 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_491 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_490 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_489 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_488 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_487 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_486 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_485 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_484 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_483 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_482 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_481 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_480 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_479 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_478 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_477 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_476 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_475 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_474 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_473 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_472 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_471 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_470 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_469 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_468 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_467 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_466 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_465 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_464 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_463 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_462 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_461 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_460 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_459 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_458 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_457 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_456 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_455 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_454 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_453 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_452 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_451 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_450 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_449 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_448 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_447 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_446 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_445 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_444 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_443 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_442 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_441 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_440 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_439 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_438 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_437 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_436 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_435 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_434 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_433 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_432 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_431 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_430 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_429 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_428 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_427 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_426 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_425 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_424 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_423 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_422 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_421 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_420 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_419 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_418 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_417 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_416 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_415 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_414 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_413 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_412 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_411 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_410 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_409 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_408 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_407 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_406 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_405 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_404 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_403 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_402 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_401 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_400 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_399 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_398 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_397 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_396 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_395 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_394 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_393 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_392 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_391 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_390 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_389 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_388 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_387 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_386 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_385 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_384 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_383 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_382 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_381 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_380 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_379 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_378 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_377 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_376 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_375 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_374 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_373 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_372 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_371 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_370 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_369 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_368 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_367 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_366 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_365 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_364 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_363 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_362 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_361 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_360 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_359 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_358 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_357 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_356 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_355 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_354 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_353 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_352 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_351 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_350 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_349 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_348 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_347 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_346 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_345 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_344 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_343 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_342 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_341 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_340 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_339 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_338 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_337 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_336 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_335 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_334 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_333 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_332 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_331 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_330 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_329 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_328 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_327 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_326 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_325 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_324 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_323 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_322 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_321 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_320 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_319 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_318 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_317 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_316 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_315 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_314 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_313 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_312 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_311 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_310 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_309 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_308 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_307 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_306 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_305 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_304 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_303 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_302 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_301 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_300 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_299 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_298 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_297 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_296 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_295 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_294 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_293 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_292 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_291 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_290 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_289 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_288 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_287 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_286 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_285 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_284 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_283 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_282 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_281 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_280 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_279 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_278 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_277 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_276 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_275 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_274 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_273 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_272 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_271 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_270 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_269 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_268 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_267 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_266 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_265 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_264 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_263 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_262 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_261 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_260 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_259 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_258 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_257 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_256 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_255 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_254 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_253 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_252 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_251 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_250 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_249 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_248 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_247 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_246 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_245 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_244 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_243 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_242 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_241 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_240 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_239 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_238 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_237 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_236 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_235 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_234 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_233 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_232 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_231 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_230 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_229 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_228 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_227 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_226 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_225 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_224 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_223 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_222 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_221 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_220 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_219 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_218 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_217 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_216 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_215 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_214 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_213 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_212 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_211 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_210 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_209 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_208 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_207 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_206 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_205 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_204 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_203 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_202 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_201 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_200 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_199 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_198 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_197 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_196 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_195 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_194 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_193 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_192 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_191 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_190 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_189 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_188 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_187 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_186 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_185 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_184 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_183 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_182 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_181 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_180 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_179 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_178 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_177 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_176 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_175 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_174 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_173 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_172 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_171 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_170 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_169 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_168 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_167 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_166 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_165 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_164 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_163 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_162 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_161 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_160 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_159 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_158 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_157 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_156 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_155 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_154 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_153 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_152 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_151 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_150 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_149 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_148 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_147 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_146 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_145 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_144 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_143 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_142 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_141 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_140 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_139 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_138 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_137 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_136 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_135 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_134 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_133 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_132 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_131 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_130 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_129 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_128 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_127 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_126 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_125 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_124 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_123 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_122 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_121 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_120 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_119 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_118 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_117 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_116 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_115 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_114 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_113 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_112 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_111 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_110 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_109 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_108 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_107 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_106 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_105 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_104 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_103 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_102 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_101 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_100 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_99 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_98 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_97 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_96 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_95 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_94 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_93 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_92 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_91 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_90 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_89 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_88 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_87 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_86 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_85 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_84 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_83 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_82 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_81 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_80 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_79 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_78 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_77 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_76 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_75 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_74 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_73 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_72 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_71 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_70 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_69 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_68 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_67 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_66 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_65 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_64 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_63 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_62 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_61 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_60 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_59 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_58 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_57 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_56 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_55 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_54 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_53 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_52 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_51 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_50 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_49 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_48 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_47 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_46 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_45 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_44 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_43 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_42 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_41 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_40 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_39 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_38 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_37 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_36 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_35 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_34 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_33 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_32 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_31 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_30 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_29 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_28 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_27 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_26 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_25 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_24 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_23 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_22 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_21 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_20 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_19 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_18 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_17 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_16 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_15 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_14 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_13 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_12 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_11 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_10 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_9 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_8 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_7 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_6 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_5 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_4 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_3 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_2 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module and_2_1 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module fa_2_159 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_350 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_349 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1373 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1372 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_675 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_158 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_348 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_347 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1371 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1370 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_674 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_157 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_346 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_345 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1369 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1368 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_673 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_156 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_344 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_343 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1367 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1366 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_672 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_155 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_342 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_341 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1365 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1364 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_671 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_154 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_340 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_339 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1363 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1362 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_670 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_153 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_338 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_337 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1361 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1360 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_669 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_152 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_336 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_335 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1359 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1358 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_668 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_151 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_334 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_333 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1357 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1356 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_667 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_150 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_332 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_331 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1355 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1354 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_666 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_149 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_330 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_329 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1353 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1352 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_665 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_148 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_328 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_327 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1351 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1350 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_664 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_147 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_326 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_325 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1349 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1348 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_663 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_146 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_324 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_323 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1347 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1346 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_662 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_145 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_322 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_321 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1345 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1344 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_661 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_144 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_320 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_319 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1343 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1342 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_660 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_143 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_318 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_317 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1341 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1340 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_659 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_142 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_316 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_315 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1339 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1338 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_658 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_141 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_314 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_313 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1337 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1336 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_657 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_140 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_312 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_311 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1335 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1334 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_656 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_139 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_310 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_309 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1333 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1332 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_655 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_138 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_308 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_307 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1331 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1330 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_654 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_137 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_306 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_305 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1329 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1328 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_653 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_136 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_304 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_303 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1327 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1326 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_652 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_135 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_302 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_301 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1325 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1324 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_651 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_134 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_300 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_299 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1323 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1322 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_650 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_133 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_298 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_297 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1321 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1320 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_649 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_132 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_296 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_295 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1319 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1318 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_648 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_131 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_294 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_293 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1317 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1316 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_647 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_130 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_292 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_291 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1315 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1314 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_646 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_129 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_290 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_289 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1313 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1312 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_645 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_128 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_288 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_287 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_352 and1 ( .a(a), .b(b), .y(s3) );
  and_2_351 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_160 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_127 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_286 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_285 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_350 and1 ( .a(a), .b(b), .y(s3) );
  and_2_349 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_159 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_126 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_284 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_283 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_348 and1 ( .a(a), .b(b), .y(s3) );
  and_2_347 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_158 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_125 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_282 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_281 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_346 and1 ( .a(a), .b(b), .y(s3) );
  and_2_345 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_157 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_124 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_280 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_279 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_344 and1 ( .a(a), .b(b), .y(s3) );
  and_2_343 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_156 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_123 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_278 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_277 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_342 and1 ( .a(a), .b(b), .y(s3) );
  and_2_341 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_155 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_122 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_276 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_275 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_340 and1 ( .a(a), .b(b), .y(s3) );
  and_2_339 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_154 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_121 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_274 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_273 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_338 and1 ( .a(a), .b(b), .y(s3) );
  and_2_337 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_153 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_120 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_272 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_271 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_336 and1 ( .a(a), .b(b), .y(s3) );
  and_2_335 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_152 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_119 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_270 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_269 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_334 and1 ( .a(a), .b(b), .y(s3) );
  and_2_333 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_151 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_118 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_268 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_267 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_332 and1 ( .a(a), .b(b), .y(s3) );
  and_2_331 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_150 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_117 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_266 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_265 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_330 and1 ( .a(a), .b(b), .y(s3) );
  and_2_329 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_149 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_116 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_264 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_263 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_328 and1 ( .a(a), .b(b), .y(s3) );
  and_2_327 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_148 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_115 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_262 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_261 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_326 and1 ( .a(a), .b(b), .y(s3) );
  and_2_325 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_147 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_114 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_260 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_259 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_324 and1 ( .a(a), .b(b), .y(s3) );
  and_2_323 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_146 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_113 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_258 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_257 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_322 and1 ( .a(a), .b(b), .y(s3) );
  and_2_321 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_145 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_112 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_256 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_255 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_320 and1 ( .a(a), .b(b), .y(s3) );
  and_2_319 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_144 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_111 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_254 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_253 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_318 and1 ( .a(a), .b(b), .y(s3) );
  and_2_317 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_143 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_110 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_252 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_251 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_316 and1 ( .a(a), .b(b), .y(s3) );
  and_2_315 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_142 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_109 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_250 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_249 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_314 and1 ( .a(a), .b(b), .y(s3) );
  and_2_313 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_141 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_108 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_248 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_247 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_312 and1 ( .a(a), .b(b), .y(s3) );
  and_2_311 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_140 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_107 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_246 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_245 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_310 and1 ( .a(a), .b(b), .y(s3) );
  and_2_309 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_139 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_106 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_244 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_243 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_308 and1 ( .a(a), .b(b), .y(s3) );
  and_2_307 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_138 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_105 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_242 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_241 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_306 and1 ( .a(a), .b(b), .y(s3) );
  and_2_305 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_137 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_104 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_240 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_239 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_304 and1 ( .a(a), .b(b), .y(s3) );
  and_2_303 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_136 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_103 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_238 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_237 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_302 and1 ( .a(a), .b(b), .y(s3) );
  and_2_301 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_135 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_102 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_236 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_235 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_300 and1 ( .a(a), .b(b), .y(s3) );
  and_2_299 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_134 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_101 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_234 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_233 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_298 and1 ( .a(a), .b(b), .y(s3) );
  and_2_297 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_133 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_100 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_232 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_231 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_296 and1 ( .a(a), .b(b), .y(s3) );
  and_2_295 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_132 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_99 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_230 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_229 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_294 and1 ( .a(a), .b(b), .y(s3) );
  and_2_293 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_131 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_98 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_228 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_227 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_292 and1 ( .a(a), .b(b), .y(s3) );
  and_2_291 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_130 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_97 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_226 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_225 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_290 and1 ( .a(a), .b(b), .y(s3) );
  and_2_289 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_129 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_96 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_224 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_223 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_288 and1 ( .a(a), .b(b), .y(s3) );
  and_2_287 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_128 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_95 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_222 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_221 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_286 and1 ( .a(a), .b(b), .y(s3) );
  and_2_285 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_127 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_94 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_220 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_219 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_284 and1 ( .a(a), .b(b), .y(s3) );
  and_2_283 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_126 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_93 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_218 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_217 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_282 and1 ( .a(a), .b(b), .y(s3) );
  and_2_281 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_125 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_92 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_216 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_215 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_280 and1 ( .a(a), .b(b), .y(s3) );
  and_2_279 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_124 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_91 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_214 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_213 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_278 and1 ( .a(a), .b(b), .y(s3) );
  and_2_277 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_123 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_90 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_212 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_211 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_276 and1 ( .a(a), .b(b), .y(s3) );
  and_2_275 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_122 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_89 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_210 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_209 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_274 and1 ( .a(a), .b(b), .y(s3) );
  and_2_273 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_121 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_88 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_208 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_207 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_272 and1 ( .a(a), .b(b), .y(s3) );
  and_2_271 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_120 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_87 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_206 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_205 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_270 and1 ( .a(a), .b(b), .y(s3) );
  and_2_269 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_119 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_86 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_204 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_203 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_268 and1 ( .a(a), .b(b), .y(s3) );
  and_2_267 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_118 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_85 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_202 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_201 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_266 and1 ( .a(a), .b(b), .y(s3) );
  and_2_265 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_117 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_84 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_200 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_199 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_264 and1 ( .a(a), .b(b), .y(s3) );
  and_2_263 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_116 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_83 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_198 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_197 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_262 and1 ( .a(a), .b(b), .y(s3) );
  and_2_261 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_115 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_82 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_196 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_195 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_260 and1 ( .a(a), .b(b), .y(s3) );
  and_2_259 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_114 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_81 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_194 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_193 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_258 and1 ( .a(a), .b(b), .y(s3) );
  and_2_257 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_113 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_80 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_192 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_191 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_256 and1 ( .a(a), .b(b), .y(s3) );
  and_2_255 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_112 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_79 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_190 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_189 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_254 and1 ( .a(a), .b(b), .y(s3) );
  and_2_253 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_111 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_78 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_188 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_187 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_252 and1 ( .a(a), .b(b), .y(s3) );
  and_2_251 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_110 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_77 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_186 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_185 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_250 and1 ( .a(a), .b(b), .y(s3) );
  and_2_249 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_109 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_76 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_184 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_183 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_248 and1 ( .a(a), .b(b), .y(s3) );
  and_2_247 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_108 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_75 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_182 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_181 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_246 and1 ( .a(a), .b(b), .y(s3) );
  and_2_245 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_107 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_74 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_180 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_179 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_244 and1 ( .a(a), .b(b), .y(s3) );
  and_2_243 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_106 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_73 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_178 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_177 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_242 and1 ( .a(a), .b(b), .y(s3) );
  and_2_241 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_105 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_72 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_176 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_175 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_240 and1 ( .a(a), .b(b), .y(s3) );
  and_2_239 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_104 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_71 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_174 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_173 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_238 and1 ( .a(a), .b(b), .y(s3) );
  and_2_237 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_103 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_70 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_172 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_171 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_236 and1 ( .a(a), .b(b), .y(s3) );
  and_2_235 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_102 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_69 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_170 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_169 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_234 and1 ( .a(a), .b(b), .y(s3) );
  and_2_233 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_101 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_68 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_168 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_167 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_232 and1 ( .a(a), .b(b), .y(s3) );
  and_2_231 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_100 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_67 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_166 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_165 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_230 and1 ( .a(a), .b(b), .y(s3) );
  and_2_229 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_99 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_66 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_164 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_163 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_228 and1 ( .a(a), .b(b), .y(s3) );
  and_2_227 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_98 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_65 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_162 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_161 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_226 and1 ( .a(a), .b(b), .y(s3) );
  and_2_225 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_97 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_64 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_128 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_127 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_192 and1 ( .a(a), .b(b), .y(s3) );
  and_2_191 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_96 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_63 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_126 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_125 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_190 and1 ( .a(a), .b(b), .y(s3) );
  and_2_189 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_95 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_62 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_124 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_123 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_188 and1 ( .a(a), .b(b), .y(s3) );
  and_2_187 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_94 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_61 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_122 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_121 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_186 and1 ( .a(a), .b(b), .y(s3) );
  and_2_185 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_93 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_60 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_120 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_119 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_184 and1 ( .a(a), .b(b), .y(s3) );
  and_2_183 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_92 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_59 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_118 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_117 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_182 and1 ( .a(a), .b(b), .y(s3) );
  and_2_181 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_91 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_58 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_116 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_115 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_180 and1 ( .a(a), .b(b), .y(s3) );
  and_2_179 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_90 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_57 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_114 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_113 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_178 and1 ( .a(a), .b(b), .y(s3) );
  and_2_177 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_89 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_56 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_112 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_111 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_168 and1 ( .a(a), .b(b), .y(s3) );
  and_2_167 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_84 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_55 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_110 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_109 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_166 and1 ( .a(a), .b(b), .y(s3) );
  and_2_165 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_83 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_54 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_108 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_107 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_164 and1 ( .a(a), .b(b), .y(s3) );
  and_2_163 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_82 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_53 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_106 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_105 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_162 and1 ( .a(a), .b(b), .y(s3) );
  and_2_161 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_81 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_52 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_104 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_103 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_160 and1 ( .a(a), .b(b), .y(s3) );
  and_2_159 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_80 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_51 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_102 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_101 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_158 and1 ( .a(a), .b(b), .y(s3) );
  and_2_157 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_79 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_50 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_100 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_99 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_156 and1 ( .a(a), .b(b), .y(s3) );
  and_2_155 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_78 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_49 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_98 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_97 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_154 and1 ( .a(a), .b(b), .y(s3) );
  and_2_153 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_77 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_48 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_96 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_95 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_144 and1 ( .a(a), .b(b), .y(s3) );
  and_2_143 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_72 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_47 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_94 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_93 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_142 and1 ( .a(a), .b(b), .y(s3) );
  and_2_141 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_71 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_46 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_92 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_91 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_140 and1 ( .a(a), .b(b), .y(s3) );
  and_2_139 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_70 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_45 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_90 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_89 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_138 and1 ( .a(a), .b(b), .y(s3) );
  and_2_137 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_69 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_44 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_88 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_87 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_136 and1 ( .a(a), .b(b), .y(s3) );
  and_2_135 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_68 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_43 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_86 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_85 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_134 and1 ( .a(a), .b(b), .y(s3) );
  and_2_133 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_67 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_42 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_84 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_83 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_132 and1 ( .a(a), .b(b), .y(s3) );
  and_2_131 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_66 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_41 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_82 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_81 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_130 and1 ( .a(a), .b(b), .y(s3) );
  and_2_129 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_65 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_40 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_80 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_79 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_120 and1 ( .a(a), .b(b), .y(s3) );
  and_2_119 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_60 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_39 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_78 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_77 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_118 and1 ( .a(a), .b(b), .y(s3) );
  and_2_117 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_59 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_38 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_76 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_75 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_116 and1 ( .a(a), .b(b), .y(s3) );
  and_2_115 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_58 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_37 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_74 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_73 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_114 and1 ( .a(a), .b(b), .y(s3) );
  and_2_113 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_57 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_36 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_72 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_71 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_112 and1 ( .a(a), .b(b), .y(s3) );
  and_2_111 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_56 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_35 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_70 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_69 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_110 and1 ( .a(a), .b(b), .y(s3) );
  and_2_109 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_55 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_34 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_68 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_67 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_108 and1 ( .a(a), .b(b), .y(s3) );
  and_2_107 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_54 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_33 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_66 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_65 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_106 and1 ( .a(a), .b(b), .y(s3) );
  and_2_105 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_53 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_32 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_64 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_63 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_96 and1 ( .a(a), .b(b), .y(s3) );
  and_2_95 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_48 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_31 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_62 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_61 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_94 and1 ( .a(a), .b(b), .y(s3) );
  and_2_93 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_47 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_30 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_60 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_59 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_92 and1 ( .a(a), .b(b), .y(s3) );
  and_2_91 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_46 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_29 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_58 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_57 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_90 and1 ( .a(a), .b(b), .y(s3) );
  and_2_89 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_45 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_28 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_56 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_55 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_88 and1 ( .a(a), .b(b), .y(s3) );
  and_2_87 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_44 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_27 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_54 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_53 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_86 and1 ( .a(a), .b(b), .y(s3) );
  and_2_85 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_43 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_26 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_52 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_51 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_84 and1 ( .a(a), .b(b), .y(s3) );
  and_2_83 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_42 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_25 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_50 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_49 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_82 and1 ( .a(a), .b(b), .y(s3) );
  and_2_81 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_41 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_24 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_48 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_47 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_72 and1 ( .a(a), .b(b), .y(s3) );
  and_2_71 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_36 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_23 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_46 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_45 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_70 and1 ( .a(a), .b(b), .y(s3) );
  and_2_69 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_35 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_22 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_44 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_43 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_68 and1 ( .a(a), .b(b), .y(s3) );
  and_2_67 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_34 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_21 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_42 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_41 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_66 and1 ( .a(a), .b(b), .y(s3) );
  and_2_65 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_33 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_20 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_40 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_39 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_64 and1 ( .a(a), .b(b), .y(s3) );
  and_2_63 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_32 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_19 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_38 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_37 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_62 and1 ( .a(a), .b(b), .y(s3) );
  and_2_61 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_31 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_18 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_36 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_35 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_60 and1 ( .a(a), .b(b), .y(s3) );
  and_2_59 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_30 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_17 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_34 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_33 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_58 and1 ( .a(a), .b(b), .y(s3) );
  and_2_57 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_29 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_16 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_32 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_31 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_48 and1 ( .a(a), .b(b), .y(s3) );
  and_2_47 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_24 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_15 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_30 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_29 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_46 and1 ( .a(a), .b(b), .y(s3) );
  and_2_45 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_23 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_14 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_28 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_27 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_44 and1 ( .a(a), .b(b), .y(s3) );
  and_2_43 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_22 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_13 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_26 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_25 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_42 and1 ( .a(a), .b(b), .y(s3) );
  and_2_41 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_21 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_12 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_24 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_23 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_40 and1 ( .a(a), .b(b), .y(s3) );
  and_2_39 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_20 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_11 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_22 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_21 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_38 and1 ( .a(a), .b(b), .y(s3) );
  and_2_37 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_19 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_10 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_20 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_19 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_36 and1 ( .a(a), .b(b), .y(s3) );
  and_2_35 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_18 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_9 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_18 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_17 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_34 and1 ( .a(a), .b(b), .y(s3) );
  and_2_33 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_17 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_8 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_16 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_15 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_24 and1 ( .a(a), .b(b), .y(s3) );
  and_2_23 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_12 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_7 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_14 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_13 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_22 and1 ( .a(a), .b(b), .y(s3) );
  and_2_21 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_11 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_6 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_12 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_11 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_20 and1 ( .a(a), .b(b), .y(s3) );
  and_2_19 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_10 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_5 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_10 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_9 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_18 and1 ( .a(a), .b(b), .y(s3) );
  and_2_17 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_9 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_4 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_8 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_7 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_16 and1 ( .a(a), .b(b), .y(s3) );
  and_2_15 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_8 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_3 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_6 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_5 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_14 and1 ( .a(a), .b(b), .y(s3) );
  and_2_13 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_7 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_2 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_4 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_3 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_12 and1 ( .a(a), .b(b), .y(s3) );
  and_2_11 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_6 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module fa_2_1 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_2 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_1 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_10 and1 ( .a(a), .b(b), .y(s3) );
  and_2_9 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_5 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module xor_2_352 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_351 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_350 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_349 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_348 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_347 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_346 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_345 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_344 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_343 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_342 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_341 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_340 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_339 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_338 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_337 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_336 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_335 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_334 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_333 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_332 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_331 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_330 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_329 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_328 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_327 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_326 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_325 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_324 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_323 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_322 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_321 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_320 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_319 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_318 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_317 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_316 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_315 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_314 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_313 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_312 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_311 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_310 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_309 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_308 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_307 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_306 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_305 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_304 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_303 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_302 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_301 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_300 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_299 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_298 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_297 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_296 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_295 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_294 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_293 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_292 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_291 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_290 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_289 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_288 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_287 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_286 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_285 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_284 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_283 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_282 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_281 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_280 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_279 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_278 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_277 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_276 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_275 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_274 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_273 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_272 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_271 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_270 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_269 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_268 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_267 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_266 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_265 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_264 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_263 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_262 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_261 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_260 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_259 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_258 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_257 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_256 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_255 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_254 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_253 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_252 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_251 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_250 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_249 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_248 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_247 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_246 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_245 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_244 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_243 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_242 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_241 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_240 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_239 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_238 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_237 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_236 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_235 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_234 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_233 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_232 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_231 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_230 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_229 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_228 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_227 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_226 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_225 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_224 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_223 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_222 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_221 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_220 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_219 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_218 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_217 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_216 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_215 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_214 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_213 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_212 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_211 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_210 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_209 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_208 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_207 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_206 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_205 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_204 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_203 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_202 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_201 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_200 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_199 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_198 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_197 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_196 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_195 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_194 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_193 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_192 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_191 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_190 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_189 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_188 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_187 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_186 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_185 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_184 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_183 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_182 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_181 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_180 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_179 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_178 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_177 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_176 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_175 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_174 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_173 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_172 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_171 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_170 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_169 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_168 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_167 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_166 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_165 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_164 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_163 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_162 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_161 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_160 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_159 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_158 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_157 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_156 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_155 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_154 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_153 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_152 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_151 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_150 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_149 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_148 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_147 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_146 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_145 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_144 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_143 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_142 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_141 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_140 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_139 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_138 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_137 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_136 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_135 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_134 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_133 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_132 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_131 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_130 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_129 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_128 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_127 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_126 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_125 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_124 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_123 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_122 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_121 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_120 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_119 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_118 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_117 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_116 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_115 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_114 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_113 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_112 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_111 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_110 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_109 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_108 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_107 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_106 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_105 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_104 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_103 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_102 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_101 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_100 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_99 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_98 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_97 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_96 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_95 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_94 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_93 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_92 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_91 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_90 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_89 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_88 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_87 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_86 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_85 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_84 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_83 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_82 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_81 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_80 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_79 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_78 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_77 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_76 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_75 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_74 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_73 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_72 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_71 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_70 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_69 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_68 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_67 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_66 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_65 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_64 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_63 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_62 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_61 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_60 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_59 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_58 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_57 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_56 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_55 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_54 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_53 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_52 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_51 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_50 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_49 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_48 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_47 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_46 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_45 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_44 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_43 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_42 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_41 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_40 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_39 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_38 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_37 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_36 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_35 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_34 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_33 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_32 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_31 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_30 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_29 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_28 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_27 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_26 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_25 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_24 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_23 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_22 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_21 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_20 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_19 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_18 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_17 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_16 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_15 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_14 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_13 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_12 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_11 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_10 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_9 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_8 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_7 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_6 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_5 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_4 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_3 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_2 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module xor_2_1 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module reg_n_n5_2 ( clock, reset, enable, x, y );
  input [4:0] x;
  output [4:0] y;
  input clock, reset, enable;


  ffd_async_74 ff_0 ( .clk(clock), .reset(reset), .en(enable), .d(x[0]), .q(
        y[0]) );
  ffd_async_73 ff_1 ( .clk(clock), .reset(reset), .en(enable), .d(x[1]), .q(
        y[1]) );
  ffd_async_72 ff_2 ( .clk(clock), .reset(reset), .en(enable), .d(x[2]), .q(
        y[2]) );
  ffd_async_71 ff_3 ( .clk(clock), .reset(reset), .en(enable), .d(x[3]), .q(
        y[3]) );
  ffd_async_70 ff_4 ( .clk(clock), .reset(reset), .en(enable), .d(x[4]), .q(
        y[4]) );
endmodule


module reg_n_n5_1 ( clock, reset, enable, x, y );
  input [4:0] x;
  output [4:0] y;
  input clock, reset, enable;


  ffd_async_5 ff_0 ( .clk(clock), .reset(reset), .en(enable), .d(x[0]), .q(
        y[0]) );
  ffd_async_4 ff_1 ( .clk(clock), .reset(reset), .en(enable), .d(x[1]), .q(
        y[1]) );
  ffd_async_3 ff_2 ( .clk(clock), .reset(reset), .en(enable), .d(x[2]), .q(
        y[2]) );
  ffd_async_2 ff_3 ( .clk(clock), .reset(reset), .en(enable), .d(x[3]), .q(
        y[3]) );
  ffd_async_1 ff_4 ( .clk(clock), .reset(reset), .en(enable), .d(x[4]), .q(
        y[4]) );
endmodule


module rca_n_n32_2 ( a, b, c_in, sum, c_out );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input c_in;
  output c_out;

  wire   [31:1] temp;

  fa_2_128 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_127 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), 
        .c_out(temp[2]) );
  fa_2_126 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), 
        .c_out(temp[3]) );
  fa_2_125 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), 
        .c_out(temp[4]) );
  fa_2_124 fa_2_i_4 ( .a(a[4]), .b(b[4]), .c_in(temp[4]), .sum(sum[4]), 
        .c_out(temp[5]) );
  fa_2_123 fa_2_i_5 ( .a(a[5]), .b(b[5]), .c_in(temp[5]), .sum(sum[5]), 
        .c_out(temp[6]) );
  fa_2_122 fa_2_i_6 ( .a(a[6]), .b(b[6]), .c_in(temp[6]), .sum(sum[6]), 
        .c_out(temp[7]) );
  fa_2_121 fa_2_i_7 ( .a(a[7]), .b(b[7]), .c_in(temp[7]), .sum(sum[7]), 
        .c_out(temp[8]) );
  fa_2_120 fa_2_i_8 ( .a(a[8]), .b(b[8]), .c_in(temp[8]), .sum(sum[8]), 
        .c_out(temp[9]) );
  fa_2_119 fa_2_i_9 ( .a(a[9]), .b(b[9]), .c_in(temp[9]), .sum(sum[9]), 
        .c_out(temp[10]) );
  fa_2_118 fa_2_i_10 ( .a(a[10]), .b(b[10]), .c_in(temp[10]), .sum(sum[10]), 
        .c_out(temp[11]) );
  fa_2_117 fa_2_i_11 ( .a(a[11]), .b(b[11]), .c_in(temp[11]), .sum(sum[11]), 
        .c_out(temp[12]) );
  fa_2_116 fa_2_i_12 ( .a(a[12]), .b(b[12]), .c_in(temp[12]), .sum(sum[12]), 
        .c_out(temp[13]) );
  fa_2_115 fa_2_i_13 ( .a(a[13]), .b(b[13]), .c_in(temp[13]), .sum(sum[13]), 
        .c_out(temp[14]) );
  fa_2_114 fa_2_i_14 ( .a(a[14]), .b(b[14]), .c_in(temp[14]), .sum(sum[14]), 
        .c_out(temp[15]) );
  fa_2_113 fa_2_i_15 ( .a(a[15]), .b(b[15]), .c_in(temp[15]), .sum(sum[15]), 
        .c_out(temp[16]) );
  fa_2_112 fa_2_i_16 ( .a(a[16]), .b(b[16]), .c_in(temp[16]), .sum(sum[16]), 
        .c_out(temp[17]) );
  fa_2_111 fa_2_i_17 ( .a(a[17]), .b(b[17]), .c_in(temp[17]), .sum(sum[17]), 
        .c_out(temp[18]) );
  fa_2_110 fa_2_i_18 ( .a(a[18]), .b(b[18]), .c_in(temp[18]), .sum(sum[18]), 
        .c_out(temp[19]) );
  fa_2_109 fa_2_i_19 ( .a(a[19]), .b(b[19]), .c_in(temp[19]), .sum(sum[19]), 
        .c_out(temp[20]) );
  fa_2_108 fa_2_i_20 ( .a(a[20]), .b(b[20]), .c_in(temp[20]), .sum(sum[20]), 
        .c_out(temp[21]) );
  fa_2_107 fa_2_i_21 ( .a(a[21]), .b(b[21]), .c_in(temp[21]), .sum(sum[21]), 
        .c_out(temp[22]) );
  fa_2_106 fa_2_i_22 ( .a(a[22]), .b(b[22]), .c_in(temp[22]), .sum(sum[22]), 
        .c_out(temp[23]) );
  fa_2_105 fa_2_i_23 ( .a(a[23]), .b(b[23]), .c_in(temp[23]), .sum(sum[23]), 
        .c_out(temp[24]) );
  fa_2_104 fa_2_i_24 ( .a(a[24]), .b(b[24]), .c_in(temp[24]), .sum(sum[24]), 
        .c_out(temp[25]) );
  fa_2_103 fa_2_i_25 ( .a(a[25]), .b(b[25]), .c_in(temp[25]), .sum(sum[25]), 
        .c_out(temp[26]) );
  fa_2_102 fa_2_i_26 ( .a(a[26]), .b(b[26]), .c_in(temp[26]), .sum(sum[26]), 
        .c_out(temp[27]) );
  fa_2_101 fa_2_i_27 ( .a(a[27]), .b(b[27]), .c_in(temp[27]), .sum(sum[27]), 
        .c_out(temp[28]) );
  fa_2_100 fa_2_i_28 ( .a(a[28]), .b(b[28]), .c_in(temp[28]), .sum(sum[28]), 
        .c_out(temp[29]) );
  fa_2_99 fa_2_i_29 ( .a(a[29]), .b(b[29]), .c_in(temp[29]), .sum(sum[29]), 
        .c_out(temp[30]) );
  fa_2_98 fa_2_i_30 ( .a(a[30]), .b(b[30]), .c_in(temp[30]), .sum(sum[30]), 
        .c_out(temp[31]) );
  fa_2_97 fa_2_i_31 ( .a(a[31]), .b(b[31]), .c_in(temp[31]), .sum(sum[31]), 
        .c_out(c_out) );
endmodule


module rca_n_n32_1 ( a, b, c_in, sum, c_out );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input c_in;
  output c_out;

  wire   [31:1] temp;

  fa_2_96 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_95 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_94 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_93 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        temp[4]) );
  fa_2_92 fa_2_i_4 ( .a(a[4]), .b(b[4]), .c_in(temp[4]), .sum(sum[4]), .c_out(
        temp[5]) );
  fa_2_91 fa_2_i_5 ( .a(a[5]), .b(b[5]), .c_in(temp[5]), .sum(sum[5]), .c_out(
        temp[6]) );
  fa_2_90 fa_2_i_6 ( .a(a[6]), .b(b[6]), .c_in(temp[6]), .sum(sum[6]), .c_out(
        temp[7]) );
  fa_2_89 fa_2_i_7 ( .a(a[7]), .b(b[7]), .c_in(temp[7]), .sum(sum[7]), .c_out(
        temp[8]) );
  fa_2_88 fa_2_i_8 ( .a(a[8]), .b(b[8]), .c_in(temp[8]), .sum(sum[8]), .c_out(
        temp[9]) );
  fa_2_87 fa_2_i_9 ( .a(a[9]), .b(b[9]), .c_in(temp[9]), .sum(sum[9]), .c_out(
        temp[10]) );
  fa_2_86 fa_2_i_10 ( .a(a[10]), .b(b[10]), .c_in(temp[10]), .sum(sum[10]), 
        .c_out(temp[11]) );
  fa_2_85 fa_2_i_11 ( .a(a[11]), .b(b[11]), .c_in(temp[11]), .sum(sum[11]), 
        .c_out(temp[12]) );
  fa_2_84 fa_2_i_12 ( .a(a[12]), .b(b[12]), .c_in(temp[12]), .sum(sum[12]), 
        .c_out(temp[13]) );
  fa_2_83 fa_2_i_13 ( .a(a[13]), .b(b[13]), .c_in(temp[13]), .sum(sum[13]), 
        .c_out(temp[14]) );
  fa_2_82 fa_2_i_14 ( .a(a[14]), .b(b[14]), .c_in(temp[14]), .sum(sum[14]), 
        .c_out(temp[15]) );
  fa_2_81 fa_2_i_15 ( .a(a[15]), .b(b[15]), .c_in(temp[15]), .sum(sum[15]), 
        .c_out(temp[16]) );
  fa_2_80 fa_2_i_16 ( .a(a[16]), .b(b[16]), .c_in(temp[16]), .sum(sum[16]), 
        .c_out(temp[17]) );
  fa_2_79 fa_2_i_17 ( .a(a[17]), .b(b[17]), .c_in(temp[17]), .sum(sum[17]), 
        .c_out(temp[18]) );
  fa_2_78 fa_2_i_18 ( .a(a[18]), .b(b[18]), .c_in(temp[18]), .sum(sum[18]), 
        .c_out(temp[19]) );
  fa_2_77 fa_2_i_19 ( .a(a[19]), .b(b[19]), .c_in(temp[19]), .sum(sum[19]), 
        .c_out(temp[20]) );
  fa_2_76 fa_2_i_20 ( .a(a[20]), .b(b[20]), .c_in(temp[20]), .sum(sum[20]), 
        .c_out(temp[21]) );
  fa_2_75 fa_2_i_21 ( .a(a[21]), .b(b[21]), .c_in(temp[21]), .sum(sum[21]), 
        .c_out(temp[22]) );
  fa_2_74 fa_2_i_22 ( .a(a[22]), .b(b[22]), .c_in(temp[22]), .sum(sum[22]), 
        .c_out(temp[23]) );
  fa_2_73 fa_2_i_23 ( .a(a[23]), .b(b[23]), .c_in(temp[23]), .sum(sum[23]), 
        .c_out(temp[24]) );
  fa_2_72 fa_2_i_24 ( .a(a[24]), .b(b[24]), .c_in(temp[24]), .sum(sum[24]), 
        .c_out(temp[25]) );
  fa_2_71 fa_2_i_25 ( .a(a[25]), .b(b[25]), .c_in(temp[25]), .sum(sum[25]), 
        .c_out(temp[26]) );
  fa_2_70 fa_2_i_26 ( .a(a[26]), .b(b[26]), .c_in(temp[26]), .sum(sum[26]), 
        .c_out(temp[27]) );
  fa_2_69 fa_2_i_27 ( .a(a[27]), .b(b[27]), .c_in(temp[27]), .sum(sum[27]), 
        .c_out(temp[28]) );
  fa_2_68 fa_2_i_28 ( .a(a[28]), .b(b[28]), .c_in(temp[28]), .sum(sum[28]), 
        .c_out(temp[29]) );
  fa_2_67 fa_2_i_29 ( .a(a[29]), .b(b[29]), .c_in(temp[29]), .sum(sum[29]), 
        .c_out(temp[30]) );
  fa_2_66 fa_2_i_30 ( .a(a[30]), .b(b[30]), .c_in(temp[30]), .sum(sum[30]), 
        .c_out(temp[31]) );
  fa_2_65 fa_2_i_31 ( .a(a[31]), .b(b[31]), .c_in(temp[31]), .sum(sum[31]), 
        .c_out(c_out) );
endmodule


module reg_n_n32_7 ( clock, reset, enable, x, y );
  input [31:0] x;
  output [31:0] y;
  input clock, reset, enable;
  wire   n1, n2, n3;

  ffd_async_239 ff_0 ( .clk(clock), .reset(n1), .en(enable), .d(x[0]), .q(y[0]) );
  ffd_async_238 ff_1 ( .clk(clock), .reset(n1), .en(enable), .d(x[1]), .q(y[1]) );
  ffd_async_237 ff_2 ( .clk(clock), .reset(n1), .en(enable), .d(x[2]), .q(y[2]) );
  ffd_async_236 ff_3 ( .clk(clock), .reset(n1), .en(enable), .d(x[3]), .q(y[3]) );
  ffd_async_235 ff_4 ( .clk(clock), .reset(n1), .en(enable), .d(x[4]), .q(y[4]) );
  ffd_async_234 ff_5 ( .clk(clock), .reset(n1), .en(enable), .d(x[5]), .q(y[5]) );
  ffd_async_233 ff_6 ( .clk(clock), .reset(n1), .en(enable), .d(x[6]), .q(y[6]) );
  ffd_async_232 ff_7 ( .clk(clock), .reset(n1), .en(enable), .d(x[7]), .q(y[7]) );
  ffd_async_231 ff_8 ( .clk(clock), .reset(n1), .en(enable), .d(x[8]), .q(y[8]) );
  ffd_async_230 ff_9 ( .clk(clock), .reset(n1), .en(enable), .d(x[9]), .q(y[9]) );
  ffd_async_229 ff_10 ( .clk(clock), .reset(n1), .en(enable), .d(x[10]), .q(
        y[10]) );
  ffd_async_228 ff_11 ( .clk(clock), .reset(n1), .en(enable), .d(x[11]), .q(
        y[11]) );
  ffd_async_227 ff_12 ( .clk(clock), .reset(n2), .en(enable), .d(x[12]), .q(
        y[12]) );
  ffd_async_226 ff_13 ( .clk(clock), .reset(n2), .en(enable), .d(x[13]), .q(
        y[13]) );
  ffd_async_225 ff_14 ( .clk(clock), .reset(n2), .en(enable), .d(x[14]), .q(
        y[14]) );
  ffd_async_224 ff_15 ( .clk(clock), .reset(n2), .en(enable), .d(x[15]), .q(
        y[15]) );
  ffd_async_223 ff_16 ( .clk(clock), .reset(n2), .en(enable), .d(x[16]), .q(
        y[16]) );
  ffd_async_222 ff_17 ( .clk(clock), .reset(n2), .en(enable), .d(x[17]), .q(
        y[17]) );
  ffd_async_221 ff_18 ( .clk(clock), .reset(n2), .en(enable), .d(x[18]), .q(
        y[18]) );
  ffd_async_220 ff_19 ( .clk(clock), .reset(n2), .en(enable), .d(x[19]), .q(
        y[19]) );
  ffd_async_219 ff_20 ( .clk(clock), .reset(n2), .en(enable), .d(x[20]), .q(
        y[20]) );
  ffd_async_218 ff_21 ( .clk(clock), .reset(n2), .en(enable), .d(x[21]), .q(
        y[21]) );
  ffd_async_217 ff_22 ( .clk(clock), .reset(n2), .en(enable), .d(x[22]), .q(
        y[22]) );
  ffd_async_216 ff_23 ( .clk(clock), .reset(n2), .en(enable), .d(x[23]), .q(
        y[23]) );
  ffd_async_215 ff_24 ( .clk(clock), .reset(n3), .en(enable), .d(x[24]), .q(
        y[24]) );
  ffd_async_214 ff_25 ( .clk(clock), .reset(n3), .en(enable), .d(x[25]), .q(
        y[25]) );
  ffd_async_213 ff_26 ( .clk(clock), .reset(n3), .en(enable), .d(x[26]), .q(
        y[26]) );
  ffd_async_212 ff_27 ( .clk(clock), .reset(n3), .en(enable), .d(x[27]), .q(
        y[27]) );
  ffd_async_211 ff_28 ( .clk(clock), .reset(n3), .en(enable), .d(x[28]), .q(
        y[28]) );
  ffd_async_210 ff_29 ( .clk(clock), .reset(n3), .en(enable), .d(x[29]), .q(
        y[29]) );
  ffd_async_209 ff_30 ( .clk(clock), .reset(n3), .en(enable), .d(x[30]), .q(
        y[30]) );
  ffd_async_208 ff_31 ( .clk(clock), .reset(n3), .en(enable), .d(x[31]), .q(
        y[31]) );
  BUF_X1 U1 ( .A(reset), .Z(n1) );
  BUF_X1 U2 ( .A(reset), .Z(n2) );
  BUF_X1 U3 ( .A(reset), .Z(n3) );
endmodule


module reg_n_n32_6 ( clock, reset, enable, x, y );
  input [31:0] x;
  output [31:0] y;
  input clock, reset, enable;
  wire   n1, n2, n3;

  ffd_async_207 ff_0 ( .clk(clock), .reset(n1), .en(enable), .d(x[0]), .q(y[0]) );
  ffd_async_206 ff_1 ( .clk(clock), .reset(n1), .en(enable), .d(x[1]), .q(y[1]) );
  ffd_async_205 ff_2 ( .clk(clock), .reset(n1), .en(enable), .d(x[2]), .q(y[2]) );
  ffd_async_204 ff_3 ( .clk(clock), .reset(n1), .en(enable), .d(x[3]), .q(y[3]) );
  ffd_async_203 ff_4 ( .clk(clock), .reset(n1), .en(enable), .d(x[4]), .q(y[4]) );
  ffd_async_202 ff_5 ( .clk(clock), .reset(n1), .en(enable), .d(x[5]), .q(y[5]) );
  ffd_async_201 ff_6 ( .clk(clock), .reset(n1), .en(enable), .d(x[6]), .q(y[6]) );
  ffd_async_200 ff_7 ( .clk(clock), .reset(n1), .en(enable), .d(x[7]), .q(y[7]) );
  ffd_async_199 ff_8 ( .clk(clock), .reset(n1), .en(enable), .d(x[8]), .q(y[8]) );
  ffd_async_198 ff_9 ( .clk(clock), .reset(n1), .en(enable), .d(x[9]), .q(y[9]) );
  ffd_async_197 ff_10 ( .clk(clock), .reset(n1), .en(enable), .d(x[10]), .q(
        y[10]) );
  ffd_async_196 ff_11 ( .clk(clock), .reset(n1), .en(enable), .d(x[11]), .q(
        y[11]) );
  ffd_async_195 ff_12 ( .clk(clock), .reset(n2), .en(enable), .d(x[12]), .q(
        y[12]) );
  ffd_async_194 ff_13 ( .clk(clock), .reset(n2), .en(enable), .d(x[13]), .q(
        y[13]) );
  ffd_async_193 ff_14 ( .clk(clock), .reset(n2), .en(enable), .d(x[14]), .q(
        y[14]) );
  ffd_async_192 ff_15 ( .clk(clock), .reset(n2), .en(enable), .d(x[15]), .q(
        y[15]) );
  ffd_async_191 ff_16 ( .clk(clock), .reset(n2), .en(enable), .d(x[16]), .q(
        y[16]) );
  ffd_async_190 ff_17 ( .clk(clock), .reset(n2), .en(enable), .d(x[17]), .q(
        y[17]) );
  ffd_async_189 ff_18 ( .clk(clock), .reset(n2), .en(enable), .d(x[18]), .q(
        y[18]) );
  ffd_async_188 ff_19 ( .clk(clock), .reset(n2), .en(enable), .d(x[19]), .q(
        y[19]) );
  ffd_async_187 ff_20 ( .clk(clock), .reset(n2), .en(enable), .d(x[20]), .q(
        y[20]) );
  ffd_async_186 ff_21 ( .clk(clock), .reset(n2), .en(enable), .d(x[21]), .q(
        y[21]) );
  ffd_async_185 ff_22 ( .clk(clock), .reset(n2), .en(enable), .d(x[22]), .q(
        y[22]) );
  ffd_async_184 ff_23 ( .clk(clock), .reset(n2), .en(enable), .d(x[23]), .q(
        y[23]) );
  ffd_async_183 ff_24 ( .clk(clock), .reset(n3), .en(enable), .d(x[24]), .q(
        y[24]) );
  ffd_async_182 ff_25 ( .clk(clock), .reset(n3), .en(enable), .d(x[25]), .q(
        y[25]) );
  ffd_async_181 ff_26 ( .clk(clock), .reset(n3), .en(enable), .d(x[26]), .q(
        y[26]) );
  ffd_async_180 ff_27 ( .clk(clock), .reset(n3), .en(enable), .d(x[27]), .q(
        y[27]) );
  ffd_async_179 ff_28 ( .clk(clock), .reset(n3), .en(enable), .d(x[28]), .q(
        y[28]) );
  ffd_async_178 ff_29 ( .clk(clock), .reset(n3), .en(enable), .d(x[29]), .q(
        y[29]) );
  ffd_async_177 ff_30 ( .clk(clock), .reset(n3), .en(enable), .d(x[30]), .q(
        y[30]) );
  ffd_async_176 ff_31 ( .clk(clock), .reset(n3), .en(enable), .d(x[31]), .q(
        y[31]) );
  BUF_X1 U1 ( .A(reset), .Z(n1) );
  BUF_X1 U2 ( .A(reset), .Z(n2) );
  BUF_X1 U3 ( .A(reset), .Z(n3) );
endmodule


module reg_n_n32_5 ( clock, reset, enable, x, y );
  input [31:0] x;
  output [31:0] y;
  input clock, reset, enable;
  wire   n1, n2, n3;

  ffd_async_175 ff_0 ( .clk(clock), .reset(n1), .en(enable), .d(x[0]), .q(y[0]) );
  ffd_async_174 ff_1 ( .clk(clock), .reset(n1), .en(enable), .d(x[1]), .q(y[1]) );
  ffd_async_173 ff_2 ( .clk(clock), .reset(n1), .en(enable), .d(x[2]), .q(y[2]) );
  ffd_async_172 ff_3 ( .clk(clock), .reset(n1), .en(enable), .d(x[3]), .q(y[3]) );
  ffd_async_171 ff_4 ( .clk(clock), .reset(n1), .en(enable), .d(x[4]), .q(y[4]) );
  ffd_async_170 ff_5 ( .clk(clock), .reset(n1), .en(enable), .d(x[5]), .q(y[5]) );
  ffd_async_169 ff_6 ( .clk(clock), .reset(n1), .en(enable), .d(x[6]), .q(y[6]) );
  ffd_async_168 ff_7 ( .clk(clock), .reset(n1), .en(enable), .d(x[7]), .q(y[7]) );
  ffd_async_167 ff_8 ( .clk(clock), .reset(n1), .en(enable), .d(x[8]), .q(y[8]) );
  ffd_async_166 ff_9 ( .clk(clock), .reset(n1), .en(enable), .d(x[9]), .q(y[9]) );
  ffd_async_165 ff_10 ( .clk(clock), .reset(n1), .en(enable), .d(x[10]), .q(
        y[10]) );
  ffd_async_164 ff_11 ( .clk(clock), .reset(n1), .en(enable), .d(x[11]), .q(
        y[11]) );
  ffd_async_163 ff_12 ( .clk(clock), .reset(n2), .en(enable), .d(x[12]), .q(
        y[12]) );
  ffd_async_162 ff_13 ( .clk(clock), .reset(n2), .en(enable), .d(x[13]), .q(
        y[13]) );
  ffd_async_161 ff_14 ( .clk(clock), .reset(n2), .en(enable), .d(x[14]), .q(
        y[14]) );
  ffd_async_160 ff_15 ( .clk(clock), .reset(n2), .en(enable), .d(x[15]), .q(
        y[15]) );
  ffd_async_159 ff_16 ( .clk(clock), .reset(n2), .en(enable), .d(x[16]), .q(
        y[16]) );
  ffd_async_158 ff_17 ( .clk(clock), .reset(n2), .en(enable), .d(x[17]), .q(
        y[17]) );
  ffd_async_157 ff_18 ( .clk(clock), .reset(n2), .en(enable), .d(x[18]), .q(
        y[18]) );
  ffd_async_156 ff_19 ( .clk(clock), .reset(n2), .en(enable), .d(x[19]), .q(
        y[19]) );
  ffd_async_155 ff_20 ( .clk(clock), .reset(n2), .en(enable), .d(x[20]), .q(
        y[20]) );
  ffd_async_154 ff_21 ( .clk(clock), .reset(n2), .en(enable), .d(x[21]), .q(
        y[21]) );
  ffd_async_153 ff_22 ( .clk(clock), .reset(n2), .en(enable), .d(x[22]), .q(
        y[22]) );
  ffd_async_152 ff_23 ( .clk(clock), .reset(n2), .en(enable), .d(x[23]), .q(
        y[23]) );
  ffd_async_151 ff_24 ( .clk(clock), .reset(n3), .en(enable), .d(x[24]), .q(
        y[24]) );
  ffd_async_150 ff_25 ( .clk(clock), .reset(n3), .en(enable), .d(x[25]), .q(
        y[25]) );
  ffd_async_149 ff_26 ( .clk(clock), .reset(n3), .en(enable), .d(x[26]), .q(
        y[26]) );
  ffd_async_148 ff_27 ( .clk(clock), .reset(n3), .en(enable), .d(x[27]), .q(
        y[27]) );
  ffd_async_147 ff_28 ( .clk(clock), .reset(n3), .en(enable), .d(x[28]), .q(
        y[28]) );
  ffd_async_146 ff_29 ( .clk(clock), .reset(n3), .en(enable), .d(x[29]), .q(
        y[29]) );
  ffd_async_145 ff_30 ( .clk(clock), .reset(n3), .en(enable), .d(x[30]), .q(
        y[30]) );
  ffd_async_144 ff_31 ( .clk(clock), .reset(n3), .en(enable), .d(x[31]), .q(
        y[31]) );
  BUF_X1 U1 ( .A(reset), .Z(n1) );
  BUF_X1 U2 ( .A(reset), .Z(n2) );
  BUF_X1 U3 ( .A(reset), .Z(n3) );
endmodule


module reg_n_n32_4 ( clock, reset, enable, x, y );
  input [31:0] x;
  output [31:0] y;
  input clock, reset, enable;
  wire   n1, n2, n3;

  ffd_async_138 ff_0 ( .clk(clock), .reset(n1), .en(enable), .d(x[0]), .q(y[0]) );
  ffd_async_137 ff_1 ( .clk(clock), .reset(n1), .en(enable), .d(x[1]), .q(y[1]) );
  ffd_async_136 ff_2 ( .clk(clock), .reset(n1), .en(enable), .d(x[2]), .q(y[2]) );
  ffd_async_135 ff_3 ( .clk(clock), .reset(n1), .en(enable), .d(x[3]), .q(y[3]) );
  ffd_async_134 ff_4 ( .clk(clock), .reset(n1), .en(enable), .d(x[4]), .q(y[4]) );
  ffd_async_133 ff_5 ( .clk(clock), .reset(n1), .en(enable), .d(x[5]), .q(y[5]) );
  ffd_async_132 ff_6 ( .clk(clock), .reset(n1), .en(enable), .d(x[6]), .q(y[6]) );
  ffd_async_131 ff_7 ( .clk(clock), .reset(n1), .en(enable), .d(x[7]), .q(y[7]) );
  ffd_async_130 ff_8 ( .clk(clock), .reset(n1), .en(enable), .d(x[8]), .q(y[8]) );
  ffd_async_129 ff_9 ( .clk(clock), .reset(n1), .en(enable), .d(x[9]), .q(y[9]) );
  ffd_async_128 ff_10 ( .clk(clock), .reset(n1), .en(enable), .d(x[10]), .q(
        y[10]) );
  ffd_async_127 ff_11 ( .clk(clock), .reset(n1), .en(enable), .d(x[11]), .q(
        y[11]) );
  ffd_async_126 ff_12 ( .clk(clock), .reset(n2), .en(enable), .d(x[12]), .q(
        y[12]) );
  ffd_async_125 ff_13 ( .clk(clock), .reset(n2), .en(enable), .d(x[13]), .q(
        y[13]) );
  ffd_async_124 ff_14 ( .clk(clock), .reset(n2), .en(enable), .d(x[14]), .q(
        y[14]) );
  ffd_async_123 ff_15 ( .clk(clock), .reset(n2), .en(enable), .d(x[15]), .q(
        y[15]) );
  ffd_async_122 ff_16 ( .clk(clock), .reset(n2), .en(enable), .d(x[16]), .q(
        y[16]) );
  ffd_async_121 ff_17 ( .clk(clock), .reset(n2), .en(enable), .d(x[17]), .q(
        y[17]) );
  ffd_async_120 ff_18 ( .clk(clock), .reset(n2), .en(enable), .d(x[18]), .q(
        y[18]) );
  ffd_async_119 ff_19 ( .clk(clock), .reset(n2), .en(enable), .d(x[19]), .q(
        y[19]) );
  ffd_async_118 ff_20 ( .clk(clock), .reset(n2), .en(enable), .d(x[20]), .q(
        y[20]) );
  ffd_async_117 ff_21 ( .clk(clock), .reset(n2), .en(enable), .d(x[21]), .q(
        y[21]) );
  ffd_async_116 ff_22 ( .clk(clock), .reset(n2), .en(enable), .d(x[22]), .q(
        y[22]) );
  ffd_async_115 ff_23 ( .clk(clock), .reset(n2), .en(enable), .d(x[23]), .q(
        y[23]) );
  ffd_async_114 ff_24 ( .clk(clock), .reset(n3), .en(enable), .d(x[24]), .q(
        y[24]) );
  ffd_async_113 ff_25 ( .clk(clock), .reset(n3), .en(enable), .d(x[25]), .q(
        y[25]) );
  ffd_async_112 ff_26 ( .clk(clock), .reset(n3), .en(enable), .d(x[26]), .q(
        y[26]) );
  ffd_async_111 ff_27 ( .clk(clock), .reset(n3), .en(enable), .d(x[27]), .q(
        y[27]) );
  ffd_async_110 ff_28 ( .clk(clock), .reset(n3), .en(enable), .d(x[28]), .q(
        y[28]) );
  ffd_async_109 ff_29 ( .clk(clock), .reset(n3), .en(enable), .d(x[29]), .q(
        y[29]) );
  ffd_async_108 ff_30 ( .clk(clock), .reset(n3), .en(enable), .d(x[30]), .q(
        y[30]) );
  ffd_async_107 ff_31 ( .clk(clock), .reset(n3), .en(enable), .d(x[31]), .q(
        y[31]) );
  BUF_X1 U1 ( .A(reset), .Z(n1) );
  BUF_X1 U2 ( .A(reset), .Z(n2) );
  BUF_X1 U3 ( .A(reset), .Z(n3) );
endmodule


module reg_n_n32_3 ( clock, reset, enable, x, y );
  input [31:0] x;
  output [31:0] y;
  input clock, reset, enable;
  wire   n1, n2, n3;

  ffd_async_106 ff_0 ( .clk(clock), .reset(n1), .en(enable), .d(x[0]), .q(y[0]) );
  ffd_async_105 ff_1 ( .clk(clock), .reset(n1), .en(enable), .d(x[1]), .q(y[1]) );
  ffd_async_104 ff_2 ( .clk(clock), .reset(n1), .en(enable), .d(x[2]), .q(y[2]) );
  ffd_async_103 ff_3 ( .clk(clock), .reset(n1), .en(enable), .d(x[3]), .q(y[3]) );
  ffd_async_102 ff_4 ( .clk(clock), .reset(n1), .en(enable), .d(x[4]), .q(y[4]) );
  ffd_async_101 ff_5 ( .clk(clock), .reset(n1), .en(enable), .d(x[5]), .q(y[5]) );
  ffd_async_100 ff_6 ( .clk(clock), .reset(n1), .en(enable), .d(x[6]), .q(y[6]) );
  ffd_async_99 ff_7 ( .clk(clock), .reset(n1), .en(enable), .d(x[7]), .q(y[7])
         );
  ffd_async_98 ff_8 ( .clk(clock), .reset(n1), .en(enable), .d(x[8]), .q(y[8])
         );
  ffd_async_97 ff_9 ( .clk(clock), .reset(n1), .en(enable), .d(x[9]), .q(y[9])
         );
  ffd_async_96 ff_10 ( .clk(clock), .reset(n1), .en(enable), .d(x[10]), .q(
        y[10]) );
  ffd_async_95 ff_11 ( .clk(clock), .reset(n1), .en(enable), .d(x[11]), .q(
        y[11]) );
  ffd_async_94 ff_12 ( .clk(clock), .reset(n2), .en(enable), .d(x[12]), .q(
        y[12]) );
  ffd_async_93 ff_13 ( .clk(clock), .reset(n2), .en(enable), .d(x[13]), .q(
        y[13]) );
  ffd_async_92 ff_14 ( .clk(clock), .reset(n2), .en(enable), .d(x[14]), .q(
        y[14]) );
  ffd_async_91 ff_15 ( .clk(clock), .reset(n2), .en(enable), .d(x[15]), .q(
        y[15]) );
  ffd_async_90 ff_16 ( .clk(clock), .reset(n2), .en(enable), .d(x[16]), .q(
        y[16]) );
  ffd_async_89 ff_17 ( .clk(clock), .reset(n2), .en(enable), .d(x[17]), .q(
        y[17]) );
  ffd_async_88 ff_18 ( .clk(clock), .reset(n2), .en(enable), .d(x[18]), .q(
        y[18]) );
  ffd_async_87 ff_19 ( .clk(clock), .reset(n2), .en(enable), .d(x[19]), .q(
        y[19]) );
  ffd_async_86 ff_20 ( .clk(clock), .reset(n2), .en(enable), .d(x[20]), .q(
        y[20]) );
  ffd_async_85 ff_21 ( .clk(clock), .reset(n2), .en(enable), .d(x[21]), .q(
        y[21]) );
  ffd_async_84 ff_22 ( .clk(clock), .reset(n2), .en(enable), .d(x[22]), .q(
        y[22]) );
  ffd_async_83 ff_23 ( .clk(clock), .reset(n2), .en(enable), .d(x[23]), .q(
        y[23]) );
  ffd_async_82 ff_24 ( .clk(clock), .reset(n3), .en(enable), .d(x[24]), .q(
        y[24]) );
  ffd_async_81 ff_25 ( .clk(clock), .reset(n3), .en(enable), .d(x[25]), .q(
        y[25]) );
  ffd_async_80 ff_26 ( .clk(clock), .reset(n3), .en(enable), .d(x[26]), .q(
        y[26]) );
  ffd_async_79 ff_27 ( .clk(clock), .reset(n3), .en(enable), .d(x[27]), .q(
        y[27]) );
  ffd_async_78 ff_28 ( .clk(clock), .reset(n3), .en(enable), .d(x[28]), .q(
        y[28]) );
  ffd_async_77 ff_29 ( .clk(clock), .reset(n3), .en(enable), .d(x[29]), .q(
        y[29]) );
  ffd_async_76 ff_30 ( .clk(clock), .reset(n3), .en(enable), .d(x[30]), .q(
        y[30]) );
  ffd_async_75 ff_31 ( .clk(clock), .reset(n3), .en(enable), .d(x[31]), .q(
        y[31]) );
  BUF_X1 U1 ( .A(reset), .Z(n1) );
  BUF_X1 U2 ( .A(reset), .Z(n2) );
  BUF_X1 U3 ( .A(reset), .Z(n3) );
endmodule


module reg_n_n32_2 ( clock, reset, enable, x, y );
  input [31:0] x;
  output [31:0] y;
  input clock, reset, enable;
  wire   n1, n2, n3;

  ffd_async_69 ff_0 ( .clk(clock), .reset(n1), .en(enable), .d(x[0]), .q(y[0])
         );
  ffd_async_68 ff_1 ( .clk(clock), .reset(n1), .en(enable), .d(x[1]), .q(y[1])
         );
  ffd_async_67 ff_2 ( .clk(clock), .reset(n1), .en(enable), .d(x[2]), .q(y[2])
         );
  ffd_async_66 ff_3 ( .clk(clock), .reset(n1), .en(enable), .d(x[3]), .q(y[3])
         );
  ffd_async_65 ff_4 ( .clk(clock), .reset(n1), .en(enable), .d(x[4]), .q(y[4])
         );
  ffd_async_64 ff_5 ( .clk(clock), .reset(n1), .en(enable), .d(x[5]), .q(y[5])
         );
  ffd_async_63 ff_6 ( .clk(clock), .reset(n1), .en(enable), .d(x[6]), .q(y[6])
         );
  ffd_async_62 ff_7 ( .clk(clock), .reset(n1), .en(enable), .d(x[7]), .q(y[7])
         );
  ffd_async_61 ff_8 ( .clk(clock), .reset(n1), .en(enable), .d(x[8]), .q(y[8])
         );
  ffd_async_60 ff_9 ( .clk(clock), .reset(n1), .en(enable), .d(x[9]), .q(y[9])
         );
  ffd_async_59 ff_10 ( .clk(clock), .reset(n1), .en(enable), .d(x[10]), .q(
        y[10]) );
  ffd_async_58 ff_11 ( .clk(clock), .reset(n1), .en(enable), .d(x[11]), .q(
        y[11]) );
  ffd_async_57 ff_12 ( .clk(clock), .reset(n2), .en(enable), .d(x[12]), .q(
        y[12]) );
  ffd_async_56 ff_13 ( .clk(clock), .reset(n2), .en(enable), .d(x[13]), .q(
        y[13]) );
  ffd_async_55 ff_14 ( .clk(clock), .reset(n2), .en(enable), .d(x[14]), .q(
        y[14]) );
  ffd_async_54 ff_15 ( .clk(clock), .reset(n2), .en(enable), .d(x[15]), .q(
        y[15]) );
  ffd_async_53 ff_16 ( .clk(clock), .reset(n2), .en(enable), .d(x[16]), .q(
        y[16]) );
  ffd_async_52 ff_17 ( .clk(clock), .reset(n2), .en(enable), .d(x[17]), .q(
        y[17]) );
  ffd_async_51 ff_18 ( .clk(clock), .reset(n2), .en(enable), .d(x[18]), .q(
        y[18]) );
  ffd_async_50 ff_19 ( .clk(clock), .reset(n2), .en(enable), .d(x[19]), .q(
        y[19]) );
  ffd_async_49 ff_20 ( .clk(clock), .reset(n2), .en(enable), .d(x[20]), .q(
        y[20]) );
  ffd_async_48 ff_21 ( .clk(clock), .reset(n2), .en(enable), .d(x[21]), .q(
        y[21]) );
  ffd_async_47 ff_22 ( .clk(clock), .reset(n2), .en(enable), .d(x[22]), .q(
        y[22]) );
  ffd_async_46 ff_23 ( .clk(clock), .reset(n2), .en(enable), .d(x[23]), .q(
        y[23]) );
  ffd_async_45 ff_24 ( .clk(clock), .reset(n3), .en(enable), .d(x[24]), .q(
        y[24]) );
  ffd_async_44 ff_25 ( .clk(clock), .reset(n3), .en(enable), .d(x[25]), .q(
        y[25]) );
  ffd_async_43 ff_26 ( .clk(clock), .reset(n3), .en(enable), .d(x[26]), .q(
        y[26]) );
  ffd_async_42 ff_27 ( .clk(clock), .reset(n3), .en(enable), .d(x[27]), .q(
        y[27]) );
  ffd_async_41 ff_28 ( .clk(clock), .reset(n3), .en(enable), .d(x[28]), .q(
        y[28]) );
  ffd_async_40 ff_29 ( .clk(clock), .reset(n3), .en(enable), .d(x[29]), .q(
        y[29]) );
  ffd_async_39 ff_30 ( .clk(clock), .reset(n3), .en(enable), .d(x[30]), .q(
        y[30]) );
  ffd_async_38 ff_31 ( .clk(clock), .reset(n3), .en(enable), .d(x[31]), .q(
        y[31]) );
  BUF_X1 U1 ( .A(reset), .Z(n1) );
  BUF_X1 U2 ( .A(reset), .Z(n2) );
  BUF_X1 U3 ( .A(reset), .Z(n3) );
endmodule


module reg_n_n32_1 ( clock, reset, enable, x, y );
  input [31:0] x;
  output [31:0] y;
  input clock, reset, enable;
  wire   n1, n2, n3;

  ffd_async_37 ff_0 ( .clk(clock), .reset(n1), .en(enable), .d(x[0]), .q(y[0])
         );
  ffd_async_36 ff_1 ( .clk(clock), .reset(n1), .en(enable), .d(x[1]), .q(y[1])
         );
  ffd_async_35 ff_2 ( .clk(clock), .reset(n1), .en(enable), .d(x[2]), .q(y[2])
         );
  ffd_async_34 ff_3 ( .clk(clock), .reset(n1), .en(enable), .d(x[3]), .q(y[3])
         );
  ffd_async_33 ff_4 ( .clk(clock), .reset(n1), .en(enable), .d(x[4]), .q(y[4])
         );
  ffd_async_32 ff_5 ( .clk(clock), .reset(n1), .en(enable), .d(x[5]), .q(y[5])
         );
  ffd_async_31 ff_6 ( .clk(clock), .reset(n1), .en(enable), .d(x[6]), .q(y[6])
         );
  ffd_async_30 ff_7 ( .clk(clock), .reset(n1), .en(enable), .d(x[7]), .q(y[7])
         );
  ffd_async_29 ff_8 ( .clk(clock), .reset(n1), .en(enable), .d(x[8]), .q(y[8])
         );
  ffd_async_28 ff_9 ( .clk(clock), .reset(n1), .en(enable), .d(x[9]), .q(y[9])
         );
  ffd_async_27 ff_10 ( .clk(clock), .reset(n1), .en(enable), .d(x[10]), .q(
        y[10]) );
  ffd_async_26 ff_11 ( .clk(clock), .reset(n1), .en(enable), .d(x[11]), .q(
        y[11]) );
  ffd_async_25 ff_12 ( .clk(clock), .reset(n2), .en(enable), .d(x[12]), .q(
        y[12]) );
  ffd_async_24 ff_13 ( .clk(clock), .reset(n2), .en(enable), .d(x[13]), .q(
        y[13]) );
  ffd_async_23 ff_14 ( .clk(clock), .reset(n2), .en(enable), .d(x[14]), .q(
        y[14]) );
  ffd_async_22 ff_15 ( .clk(clock), .reset(n2), .en(enable), .d(x[15]), .q(
        y[15]) );
  ffd_async_21 ff_16 ( .clk(clock), .reset(n2), .en(enable), .d(x[16]), .q(
        y[16]) );
  ffd_async_20 ff_17 ( .clk(clock), .reset(n2), .en(enable), .d(x[17]), .q(
        y[17]) );
  ffd_async_19 ff_18 ( .clk(clock), .reset(n2), .en(enable), .d(x[18]), .q(
        y[18]) );
  ffd_async_18 ff_19 ( .clk(clock), .reset(n2), .en(enable), .d(x[19]), .q(
        y[19]) );
  ffd_async_17 ff_20 ( .clk(clock), .reset(n2), .en(enable), .d(x[20]), .q(
        y[20]) );
  ffd_async_16 ff_21 ( .clk(clock), .reset(n2), .en(enable), .d(x[21]), .q(
        y[21]) );
  ffd_async_15 ff_22 ( .clk(clock), .reset(n2), .en(enable), .d(x[22]), .q(
        y[22]) );
  ffd_async_14 ff_23 ( .clk(clock), .reset(n2), .en(enable), .d(x[23]), .q(
        y[23]) );
  ffd_async_13 ff_24 ( .clk(clock), .reset(n3), .en(enable), .d(x[24]), .q(
        y[24]) );
  ffd_async_12 ff_25 ( .clk(clock), .reset(n3), .en(enable), .d(x[25]), .q(
        y[25]) );
  ffd_async_11 ff_26 ( .clk(clock), .reset(n3), .en(enable), .d(x[26]), .q(
        y[26]) );
  ffd_async_10 ff_27 ( .clk(clock), .reset(n3), .en(enable), .d(x[27]), .q(
        y[27]) );
  ffd_async_9 ff_28 ( .clk(clock), .reset(n3), .en(enable), .d(x[28]), .q(
        y[28]) );
  ffd_async_8 ff_29 ( .clk(clock), .reset(n3), .en(enable), .d(x[29]), .q(
        y[29]) );
  ffd_async_7 ff_30 ( .clk(clock), .reset(n3), .en(enable), .d(x[30]), .q(
        y[30]) );
  ffd_async_6 ff_31 ( .clk(clock), .reset(n3), .en(enable), .d(x[31]), .q(
        y[31]) );
  BUF_X1 U1 ( .A(reset), .Z(n1) );
  BUF_X1 U2 ( .A(reset), .Z(n2) );
  BUF_X1 U3 ( .A(reset), .Z(n3) );
endmodule


module mux21_generic_n4_0 ( a, b, sel, y );
  input [3:0] a;
  input [3:0] b;
  output [3:0] y;
  input sel;


  mux21_32 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(sel), .y(y[0]) );
  mux21_31 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(sel), .y(y[1]) );
  mux21_30 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(sel), .y(y[2]) );
  mux21_29 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(sel), .y(y[3]) );
endmodule


module rca_n_n4_0 ( a, b, c_in, sum, c_out );
  input [3:0] a;
  input [3:0] b;
  output [3:0] sum;
  input c_in;
  output c_out;

  wire   [3:1] temp;

  fa_2_64 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_63 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), .c_out(
        temp[2]) );
  fa_2_62 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), .c_out(
        temp[3]) );
  fa_2_61 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), .c_out(
        c_out) );
endmodule


module PG_0 ( a, b, g, p );
  input a, b;
  output g, p;


  and_2_224 and_gen ( .a(a), .b(b), .y(g) );
  xor_2_160 xor_pro ( .a(a), .b(b), .y(p) );
endmodule


module carry_select_block_n4_0 ( a, b, cin, s );
  input [3:0] a;
  input [3:0] b;
  output [3:0] s;
  input cin;

  wire   [3:0] sum_first_rca;
  wire   [3:0] sum_second_rca;

  rca_n_n4_0 first_rca ( .a(a), .b(b), .c_in(1'b0), .sum(sum_first_rca) );
  rca_n_n4_15 second_rca ( .a(a), .b(b), .c_in(1'b1), .sum(sum_second_rca) );
  mux21_generic_n4_0 mux ( .a(sum_first_rca), .b(sum_second_rca), .sel(cin), 
        .y(s) );
endmodule


module PG_general_0 ( gkminj, pkminj, gik, pik, gij, pij );
  input gkminj, pkminj, gik, pik;
  output gij, pij;
  wire   and_out;

  and_2_414 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_195 or_gen ( .a(gik), .b(and_out), .y(gij) );
  and_2_413 and_prop ( .a(pik), .b(pkminj), .y(pij) );
endmodule


module G_general_0 ( gkminj, gik, pik, gij );
  input gkminj, gik, pik;
  output gij;
  wire   and_out;

  and_2_415 and_gen ( .a(pik), .b(gkminj), .y(and_out) );
  or_2_196 or_gen ( .a(gik), .b(and_out), .y(gij) );
endmodule


module PG_network_n32 ( a_n, b_n, g_n, p_n );
  input [31:0] a_n;
  input [31:0] b_n;
  output [31:0] g_n;
  output [31:0] p_n;


  PG_0 PG_i_0 ( .a(a_n[0]), .b(b_n[0]), .g(g_n[0]), .p(p_n[0]) );
  PG_31 PG_i_1 ( .a(a_n[1]), .b(b_n[1]), .g(g_n[1]), .p(p_n[1]) );
  PG_30 PG_i_2 ( .a(a_n[2]), .b(b_n[2]), .g(g_n[2]), .p(p_n[2]) );
  PG_29 PG_i_3 ( .a(a_n[3]), .b(b_n[3]), .g(g_n[3]), .p(p_n[3]) );
  PG_28 PG_i_4 ( .a(a_n[4]), .b(b_n[4]), .g(g_n[4]), .p(p_n[4]) );
  PG_27 PG_i_5 ( .a(a_n[5]), .b(b_n[5]), .g(g_n[5]), .p(p_n[5]) );
  PG_26 PG_i_6 ( .a(a_n[6]), .b(b_n[6]), .g(g_n[6]), .p(p_n[6]) );
  PG_25 PG_i_7 ( .a(a_n[7]), .b(b_n[7]), .g(g_n[7]), .p(p_n[7]) );
  PG_24 PG_i_8 ( .a(a_n[8]), .b(b_n[8]), .g(g_n[8]), .p(p_n[8]) );
  PG_23 PG_i_9 ( .a(a_n[9]), .b(b_n[9]), .g(g_n[9]), .p(p_n[9]) );
  PG_22 PG_i_10 ( .a(a_n[10]), .b(b_n[10]), .g(g_n[10]), .p(p_n[10]) );
  PG_21 PG_i_11 ( .a(a_n[11]), .b(b_n[11]), .g(g_n[11]), .p(p_n[11]) );
  PG_20 PG_i_12 ( .a(a_n[12]), .b(b_n[12]), .g(g_n[12]), .p(p_n[12]) );
  PG_19 PG_i_13 ( .a(a_n[13]), .b(b_n[13]), .g(g_n[13]), .p(p_n[13]) );
  PG_18 PG_i_14 ( .a(a_n[14]), .b(b_n[14]), .g(g_n[14]), .p(p_n[14]) );
  PG_17 PG_i_15 ( .a(a_n[15]), .b(b_n[15]), .g(g_n[15]), .p(p_n[15]) );
  PG_16 PG_i_16 ( .a(a_n[16]), .b(b_n[16]), .g(g_n[16]), .p(p_n[16]) );
  PG_15 PG_i_17 ( .a(a_n[17]), .b(b_n[17]), .g(g_n[17]), .p(p_n[17]) );
  PG_14 PG_i_18 ( .a(a_n[18]), .b(b_n[18]), .g(g_n[18]), .p(p_n[18]) );
  PG_13 PG_i_19 ( .a(a_n[19]), .b(b_n[19]), .g(g_n[19]), .p(p_n[19]) );
  PG_12 PG_i_20 ( .a(a_n[20]), .b(b_n[20]), .g(g_n[20]), .p(p_n[20]) );
  PG_11 PG_i_21 ( .a(a_n[21]), .b(b_n[21]), .g(g_n[21]), .p(p_n[21]) );
  PG_10 PG_i_22 ( .a(a_n[22]), .b(b_n[22]), .g(g_n[22]), .p(p_n[22]) );
  PG_9 PG_i_23 ( .a(a_n[23]), .b(b_n[23]), .g(g_n[23]), .p(p_n[23]) );
  PG_8 PG_i_24 ( .a(a_n[24]), .b(b_n[24]), .g(g_n[24]), .p(p_n[24]) );
  PG_7 PG_i_25 ( .a(a_n[25]), .b(b_n[25]), .g(g_n[25]), .p(p_n[25]) );
  PG_6 PG_i_26 ( .a(a_n[26]), .b(b_n[26]), .g(g_n[26]), .p(p_n[26]) );
  PG_5 PG_i_27 ( .a(a_n[27]), .b(b_n[27]), .g(g_n[27]), .p(p_n[27]) );
  PG_4 PG_i_28 ( .a(a_n[28]), .b(b_n[28]), .g(g_n[28]), .p(p_n[28]) );
  PG_3 PG_i_29 ( .a(a_n[29]), .b(b_n[29]), .g(g_n[29]), .p(p_n[29]) );
  PG_2 PG_i_30 ( .a(a_n[30]), .b(b_n[30]), .g(g_n[30]), .p(p_n[30]) );
  PG_1 PG_i_31 ( .a(a_n[31]), .b(b_n[31]), .g(g_n[31]), .p(p_n[31]) );
endmodule


module logic_0 ( r1, r2, s0, s1, s2, s3, y );
  input r1, r2, s0, s1, s2, s3;
  output y;
  wire   n3, n5, n6, n4;

  OAI22_X1 U1 ( .A1(n3), .A2(n4), .B1(r2), .B2(n5), .ZN(y) );
  AOI22_X1 U2 ( .A1(s1), .A2(n6), .B1(s3), .B2(r1), .ZN(n3) );
  AOI22_X1 U3 ( .A1(s0), .A2(n6), .B1(s2), .B2(r1), .ZN(n5) );
  INV_X1 U4 ( .A(r1), .ZN(n6) );
  INV_X1 U5 ( .A(r2), .ZN(n4) );
endmodule


module nor_n1_n32 ( a, y );
  input [31:0] a;
  output y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR4_X1 U1 ( .A1(a[5]), .A2(a[4]), .A3(a[3]), .A4(a[31]), .ZN(n9) );
  NOR4_X1 U2 ( .A1(a[30]), .A2(a[2]), .A3(a[29]), .A4(a[28]), .ZN(n8) );
  NOR4_X1 U3 ( .A1(a[23]), .A2(a[22]), .A3(a[21]), .A4(a[20]), .ZN(n6) );
  NOR4_X1 U4 ( .A1(a[27]), .A2(a[26]), .A3(a[25]), .A4(a[24]), .ZN(n7) );
  NOR4_X1 U5 ( .A1(a[9]), .A2(a[8]), .A3(a[7]), .A4(a[6]), .ZN(n10) );
  NOR4_X1 U6 ( .A1(a[16]), .A2(a[15]), .A3(a[14]), .A4(a[13]), .ZN(n4) );
  NOR2_X1 U7 ( .A1(n1), .A2(n2), .ZN(y) );
  NAND4_X1 U8 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NAND4_X1 U9 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NOR4_X1 U10 ( .A1(a[12]), .A2(a[11]), .A3(a[10]), .A4(a[0]), .ZN(n3) );
  NOR4_X1 U11 ( .A1(a[1]), .A2(a[19]), .A3(a[18]), .A4(a[17]), .ZN(n5) );
endmodule


module not_n_n32_0 ( a, y );
  input [31:0] a;
  output [31:0] y;


  not_1_416 not_1_component_0 ( .a(a[0]), .y(y[0]) );
  not_1_415 not_1_component_1 ( .a(a[1]), .y(y[1]) );
  not_1_414 not_1_component_2 ( .a(a[2]), .y(y[2]) );
  not_1_413 not_1_component_3 ( .a(a[3]), .y(y[3]) );
  not_1_412 not_1_component_4 ( .a(a[4]), .y(y[4]) );
  not_1_411 not_1_component_5 ( .a(a[5]), .y(y[5]) );
  not_1_410 not_1_component_6 ( .a(a[6]), .y(y[6]) );
  not_1_409 not_1_component_7 ( .a(a[7]), .y(y[7]) );
  not_1_408 not_1_component_8 ( .a(a[8]), .y(y[8]) );
  not_1_407 not_1_component_9 ( .a(a[9]), .y(y[9]) );
  not_1_406 not_1_component_10 ( .a(a[10]), .y(y[10]) );
  not_1_405 not_1_component_11 ( .a(a[11]), .y(y[11]) );
  not_1_404 not_1_component_12 ( .a(a[12]), .y(y[12]) );
  not_1_403 not_1_component_13 ( .a(a[13]), .y(y[13]) );
  not_1_402 not_1_component_14 ( .a(a[14]), .y(y[14]) );
  not_1_401 not_1_component_15 ( .a(a[15]), .y(y[15]) );
  not_1_400 not_1_component_16 ( .a(a[16]), .y(y[16]) );
  not_1_399 not_1_component_17 ( .a(a[17]), .y(y[17]) );
  not_1_398 not_1_component_18 ( .a(a[18]), .y(y[18]) );
  not_1_397 not_1_component_19 ( .a(a[19]), .y(y[19]) );
  not_1_396 not_1_component_20 ( .a(a[20]), .y(y[20]) );
  not_1_395 not_1_component_21 ( .a(a[21]), .y(y[21]) );
  not_1_394 not_1_component_22 ( .a(a[22]), .y(y[22]) );
  not_1_393 not_1_component_23 ( .a(a[23]), .y(y[23]) );
  not_1_392 not_1_component_24 ( .a(a[24]), .y(y[24]) );
  not_1_391 not_1_component_25 ( .a(a[25]), .y(y[25]) );
  not_1_390 not_1_component_26 ( .a(a[26]), .y(y[26]) );
  not_1_389 not_1_component_27 ( .a(a[27]), .y(y[27]) );
  not_1_388 not_1_component_28 ( .a(a[28]), .y(y[28]) );
  not_1_387 not_1_component_29 ( .a(a[29]), .y(y[29]) );
  not_1_386 not_1_component_30 ( .a(a[30]), .y(y[30]) );
  not_1_385 not_1_component_31 ( .a(a[31]), .y(y[31]) );
endmodule


module sum_generator_n32 ( a, b, c, cin, s, cout );
  input [31:0] a;
  input [31:0] b;
  input [31:0] c;
  output [31:0] s;
  input cin;
  output cout;

  assign cout = c[7];

  carry_select_block_n4_0 carry_select_block_0 ( .a(a[3:0]), .b(b[3:0]), .cin(
        cin), .s(s[3:0]) );
  carry_select_block_n4_7 carry_select_block_i_1 ( .a(a[7:4]), .b(b[7:4]), 
        .cin(c[0]), .s(s[7:4]) );
  carry_select_block_n4_6 carry_select_block_i_2 ( .a(a[11:8]), .b(b[11:8]), 
        .cin(c[1]), .s(s[11:8]) );
  carry_select_block_n4_5 carry_select_block_i_3 ( .a(a[15:12]), .b(b[15:12]), 
        .cin(c[2]), .s(s[15:12]) );
  carry_select_block_n4_4 carry_select_block_i_4 ( .a(a[19:16]), .b(b[19:16]), 
        .cin(c[3]), .s(s[19:16]) );
  carry_select_block_n4_3 carry_select_block_i_5 ( .a(a[23:20]), .b(b[23:20]), 
        .cin(c[4]), .s(s[23:20]) );
  carry_select_block_n4_2 carry_select_block_i_6 ( .a(a[27:24]), .b(b[27:24]), 
        .cin(c[5]), .s(s[27:24]) );
  carry_select_block_n4_1 carry_select_block_i_7 ( .a(a[31:28]), .b(b[31:28]), 
        .cin(c[6]), .s(s[31:28]) );
endmodule


module sparse_tree_carry_gen_n32 ( a, b, c );
  input [31:0] a;
  input [31:0] b;
  output [31:0] c;
  wire   \temp[9][7] , \temp[9][6] , \temp[8][7] , \temp[8][6] , \temp[7][7] ,
         \temp[7][5] , \temp[7][3] , \temp[6][7] , \temp[6][5] , \temp[6][3] ,
         \temp[5][7] , \temp[5][6] , \temp[5][5] , \temp[5][4] , \temp[5][3] ,
         \temp[5][2] , \temp[5][1] , \temp[4][7] , \temp[4][6] , \temp[4][5] ,
         \temp[4][4] , \temp[4][3] , \temp[4][2] , \temp[4][1] , \temp[3][15] ,
         \temp[3][14] , \temp[3][13] , \temp[3][12] , \temp[3][11] ,
         \temp[3][10] , \temp[3][9] , \temp[3][8] , \temp[3][7] , \temp[3][6] ,
         \temp[3][5] , \temp[3][4] , \temp[3][3] , \temp[3][2] , \temp[3][1] ,
         \temp[2][15] , \temp[2][14] , \temp[2][13] , \temp[2][12] ,
         \temp[2][11] , \temp[2][10] , \temp[2][9] , \temp[2][8] ,
         \temp[2][7] , \temp[2][6] , \temp[2][5] , \temp[2][4] , \temp[2][3] ,
         \temp[2][2] , \temp[2][1] , \temp[2][0] , \temp[1][31] ,
         \temp[1][30] , \temp[1][29] , \temp[1][28] , \temp[1][27] ,
         \temp[1][26] , \temp[1][25] , \temp[1][24] , \temp[1][23] ,
         \temp[1][22] , \temp[1][21] , \temp[1][20] , \temp[1][19] ,
         \temp[1][18] , \temp[1][17] , \temp[1][16] , \temp[1][15] ,
         \temp[1][14] , \temp[1][13] , \temp[1][12] , \temp[1][11] ,
         \temp[1][10] , \temp[1][9] , \temp[1][8] , \temp[1][7] , \temp[1][6] ,
         \temp[1][5] , \temp[1][4] , \temp[1][3] , \temp[1][2] , \temp[1][1] ,
         \temp[0][31] , \temp[0][30] , \temp[0][29] , \temp[0][28] ,
         \temp[0][27] , \temp[0][26] , \temp[0][25] , \temp[0][24] ,
         \temp[0][23] , \temp[0][22] , \temp[0][21] , \temp[0][20] ,
         \temp[0][19] , \temp[0][18] , \temp[0][17] , \temp[0][16] ,
         \temp[0][15] , \temp[0][14] , \temp[0][13] , \temp[0][12] ,
         \temp[0][11] , \temp[0][10] , \temp[0][9] , \temp[0][8] ,
         \temp[0][7] , \temp[0][6] , \temp[0][5] , \temp[0][4] , \temp[0][3] ,
         \temp[0][2] , \temp[0][1] , \temp[0][0] ;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign c[8] = 1'b0;
  assign c[9] = 1'b0;
  assign c[10] = 1'b0;
  assign c[11] = 1'b0;
  assign c[12] = 1'b0;
  assign c[13] = 1'b0;
  assign c[14] = 1'b0;
  assign c[15] = 1'b0;
  assign c[16] = 1'b0;
  assign c[17] = 1'b0;
  assign c[18] = 1'b0;
  assign c[19] = 1'b0;
  assign c[20] = 1'b0;
  assign c[21] = 1'b0;
  assign c[22] = 1'b0;
  assign c[23] = 1'b0;
  assign c[24] = 1'b0;
  assign c[25] = 1'b0;
  assign c[26] = 1'b0;
  assign c[27] = 1'b0;
  assign c[28] = 1'b0;
  assign c[29] = 1'b0;
  assign c[30] = 1'b0;
  assign c[31] = 1'b0;

  PG_network_n32 pg_net ( .a_n(a), .b_n(b), .g_n({\temp[0][31] , \temp[0][30] , 
        \temp[0][29] , \temp[0][28] , \temp[0][27] , \temp[0][26] , 
        \temp[0][25] , \temp[0][24] , \temp[0][23] , \temp[0][22] , 
        \temp[0][21] , \temp[0][20] , \temp[0][19] , \temp[0][18] , 
        \temp[0][17] , \temp[0][16] , \temp[0][15] , \temp[0][14] , 
        \temp[0][13] , \temp[0][12] , \temp[0][11] , \temp[0][10] , 
        \temp[0][9] , \temp[0][8] , \temp[0][7] , \temp[0][6] , \temp[0][5] , 
        \temp[0][4] , \temp[0][3] , \temp[0][2] , \temp[0][1] , \temp[0][0] }), 
        .p_n({\temp[1][31] , \temp[1][30] , \temp[1][29] , \temp[1][28] , 
        \temp[1][27] , \temp[1][26] , \temp[1][25] , \temp[1][24] , 
        \temp[1][23] , \temp[1][22] , \temp[1][21] , \temp[1][20] , 
        \temp[1][19] , \temp[1][18] , \temp[1][17] , \temp[1][16] , 
        \temp[1][15] , \temp[1][14] , \temp[1][13] , \temp[1][12] , 
        \temp[1][11] , \temp[1][10] , \temp[1][9] , \temp[1][8] , \temp[1][7] , 
        \temp[1][6] , \temp[1][5] , \temp[1][4] , \temp[1][3] , \temp[1][2] , 
        \temp[1][1] , SYNOPSYS_UNCONNECTED__0}) );
  G_general_0 gen_in_i_0 ( .gkminj(\temp[0][0] ), .gik(\temp[0][1] ), .pik(
        \temp[1][1] ), .gij(\temp[2][0] ) );
  PG_general_0 pg_j_0_0 ( .gkminj(\temp[0][2] ), .pkminj(\temp[1][2] ), .gik(
        \temp[0][3] ), .pik(\temp[1][3] ), .gij(\temp[2][1] ), .pij(
        \temp[3][1] ) );
  PG_general_26 pg_j_0_1 ( .gkminj(\temp[0][4] ), .pkminj(\temp[1][4] ), .gik(
        \temp[0][5] ), .pik(\temp[1][5] ), .gij(\temp[2][2] ), .pij(
        \temp[3][2] ) );
  PG_general_25 pg_j_0_2 ( .gkminj(\temp[0][6] ), .pkminj(\temp[1][6] ), .gik(
        \temp[0][7] ), .pik(\temp[1][7] ), .gij(\temp[2][3] ), .pij(
        \temp[3][3] ) );
  PG_general_24 pg_j_0_3 ( .gkminj(\temp[0][8] ), .pkminj(\temp[1][8] ), .gik(
        \temp[0][9] ), .pik(\temp[1][9] ), .gij(\temp[2][4] ), .pij(
        \temp[3][4] ) );
  PG_general_23 pg_j_0_4 ( .gkminj(\temp[0][10] ), .pkminj(\temp[1][10] ), 
        .gik(\temp[0][11] ), .pik(\temp[1][11] ), .gij(\temp[2][5] ), .pij(
        \temp[3][5] ) );
  PG_general_22 pg_j_0_5 ( .gkminj(\temp[0][12] ), .pkminj(\temp[1][12] ), 
        .gik(\temp[0][13] ), .pik(\temp[1][13] ), .gij(\temp[2][6] ), .pij(
        \temp[3][6] ) );
  PG_general_21 pg_j_0_6 ( .gkminj(\temp[0][14] ), .pkminj(\temp[1][14] ), 
        .gik(\temp[0][15] ), .pik(\temp[1][15] ), .gij(\temp[2][7] ), .pij(
        \temp[3][7] ) );
  PG_general_20 pg_j_0_7 ( .gkminj(\temp[0][16] ), .pkminj(\temp[1][16] ), 
        .gik(\temp[0][17] ), .pik(\temp[1][17] ), .gij(\temp[2][8] ), .pij(
        \temp[3][8] ) );
  PG_general_19 pg_j_0_8 ( .gkminj(\temp[0][18] ), .pkminj(\temp[1][18] ), 
        .gik(\temp[0][19] ), .pik(\temp[1][19] ), .gij(\temp[2][9] ), .pij(
        \temp[3][9] ) );
  PG_general_18 pg_j_0_9 ( .gkminj(\temp[0][20] ), .pkminj(\temp[1][20] ), 
        .gik(\temp[0][21] ), .pik(\temp[1][21] ), .gij(\temp[2][10] ), .pij(
        \temp[3][10] ) );
  PG_general_17 pg_j_0_10 ( .gkminj(\temp[0][22] ), .pkminj(\temp[1][22] ), 
        .gik(\temp[0][23] ), .pik(\temp[1][23] ), .gij(\temp[2][11] ), .pij(
        \temp[3][11] ) );
  PG_general_16 pg_j_0_11 ( .gkminj(\temp[0][24] ), .pkminj(\temp[1][24] ), 
        .gik(\temp[0][25] ), .pik(\temp[1][25] ), .gij(\temp[2][12] ), .pij(
        \temp[3][12] ) );
  PG_general_15 pg_j_0_12 ( .gkminj(\temp[0][26] ), .pkminj(\temp[1][26] ), 
        .gik(\temp[0][27] ), .pik(\temp[1][27] ), .gij(\temp[2][13] ), .pij(
        \temp[3][13] ) );
  PG_general_14 pg_j_0_13 ( .gkminj(\temp[0][28] ), .pkminj(\temp[1][28] ), 
        .gik(\temp[0][29] ), .pik(\temp[1][29] ), .gij(\temp[2][14] ), .pij(
        \temp[3][14] ) );
  PG_general_13 pg_j_0_14 ( .gkminj(\temp[0][30] ), .pkminj(\temp[1][30] ), 
        .gik(\temp[0][31] ), .pik(\temp[1][31] ), .gij(\temp[2][15] ), .pij(
        \temp[3][15] ) );
  G_general_8 gen_in_i_1 ( .gkminj(\temp[2][0] ), .gik(\temp[2][1] ), .pik(
        \temp[3][1] ), .gij(c[0]) );
  PG_general_12 pg_j_1_0 ( .gkminj(\temp[2][2] ), .pkminj(\temp[3][2] ), .gik(
        \temp[2][3] ), .pik(\temp[3][3] ), .gij(\temp[4][1] ), .pij(
        \temp[5][1] ) );
  PG_general_11 pg_j_1_1 ( .gkminj(\temp[2][4] ), .pkminj(\temp[3][4] ), .gik(
        \temp[2][5] ), .pik(\temp[3][5] ), .gij(\temp[4][2] ), .pij(
        \temp[5][2] ) );
  PG_general_10 pg_j_1_2 ( .gkminj(\temp[2][6] ), .pkminj(\temp[3][6] ), .gik(
        \temp[2][7] ), .pik(\temp[3][7] ), .gij(\temp[4][3] ), .pij(
        \temp[5][3] ) );
  PG_general_9 pg_j_1_3 ( .gkminj(\temp[2][8] ), .pkminj(\temp[3][8] ), .gik(
        \temp[2][9] ), .pik(\temp[3][9] ), .gij(\temp[4][4] ), .pij(
        \temp[5][4] ) );
  PG_general_8 pg_j_1_4 ( .gkminj(\temp[2][10] ), .pkminj(\temp[3][10] ), 
        .gik(\temp[2][11] ), .pik(\temp[3][11] ), .gij(\temp[4][5] ), .pij(
        \temp[5][5] ) );
  PG_general_7 pg_j_1_5 ( .gkminj(\temp[2][12] ), .pkminj(\temp[3][12] ), 
        .gik(\temp[2][13] ), .pik(\temp[3][13] ), .gij(\temp[4][6] ), .pij(
        \temp[5][6] ) );
  PG_general_6 pg_j_1_6 ( .gkminj(\temp[2][14] ), .pkminj(\temp[3][14] ), 
        .gik(\temp[2][15] ), .pik(\temp[3][15] ), .gij(\temp[4][7] ), .pij(
        \temp[5][7] ) );
  G_general_7 gen_r_2_0 ( .gkminj(c[0]), .gik(\temp[4][1] ), .pik(\temp[5][1] ), .gij(c[1]) );
  PG_general_5 pg_e_2_0_0 ( .gkminj(\temp[4][2] ), .pkminj(\temp[5][2] ), 
        .gik(\temp[4][3] ), .pik(\temp[5][3] ), .gij(\temp[6][3] ), .pij(
        \temp[7][3] ) );
  PG_general_4 pg_e_2_1_0 ( .gkminj(\temp[4][4] ), .pkminj(\temp[5][4] ), 
        .gik(\temp[4][5] ), .pik(\temp[5][5] ), .gij(\temp[6][5] ), .pij(
        \temp[7][5] ) );
  PG_general_3 pg_e_2_2_0 ( .gkminj(\temp[4][6] ), .pkminj(\temp[5][6] ), 
        .gik(\temp[4][7] ), .pik(\temp[5][7] ), .gij(\temp[6][7] ), .pij(
        \temp[7][7] ) );
  G_general_6 gen_r_3_0 ( .gkminj(c[1]), .gik(\temp[4][2] ), .pik(\temp[5][2] ), .gij(c[2]) );
  G_general_5 gen_r_3_1 ( .gkminj(c[1]), .gik(\temp[6][3] ), .pik(\temp[7][3] ), .gij(c[3]) );
  PG_general_2 pg_e_3_0_0 ( .gkminj(\temp[4][4] ), .pkminj(\temp[5][4] ), 
        .gik(\temp[4][6] ), .pik(\temp[5][6] ), .gij(\temp[8][6] ), .pij(
        \temp[9][6] ) );
  PG_general_1 pg_e_3_0_1 ( .gkminj(\temp[4][4] ), .pkminj(\temp[5][4] ), 
        .gik(\temp[6][7] ), .pik(\temp[7][7] ), .gij(\temp[8][7] ), .pij(
        \temp[9][7] ) );
  G_general_4 gen_r_4_0 ( .gkminj(c[3]), .gik(\temp[4][4] ), .pik(\temp[5][4] ), .gij(c[4]) );
  G_general_3 gen_r_4_1 ( .gkminj(c[3]), .gik(\temp[6][5] ), .pik(\temp[7][5] ), .gij(c[5]) );
  G_general_2 gen_r_4_2 ( .gkminj(c[3]), .gik(\temp[8][6] ), .pik(\temp[9][6] ), .gij(c[6]) );
  G_general_1 gen_r_4_3 ( .gkminj(c[3]), .gik(\temp[8][7] ), .pik(\temp[9][7] ), .gij(c[7]) );
endmodule


module not_1_0 ( a, y );
  input a;
  output y;


  INV_X1 U1 ( .A(a), .ZN(y) );
endmodule


module or_2_0 ( a, b, y );
  input a, b;
  output y;


  OR2_X1 U1 ( .A1(a), .A2(b), .ZN(y) );
endmodule


module and_2_1375 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module encoder_n32 ( out_add, out_sub, out_sl, out_sr, out_log, out_cmp, 
        out_eq, sel, o );
  input [31:0] out_add;
  input [31:0] out_sub;
  input [31:0] out_sl;
  input [31:0] out_sr;
  input [31:0] out_log;
  input [31:0] out_cmp;
  input [31:0] out_eq;
  input [3:0] sel;
  output [31:0] o;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n83, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107;
  tri   [31:0] out_sl;

  INV_X1 U2 ( .A(out_eq[0]), .ZN(n81) );
  NAND2_X1 U3 ( .A1(out_cmp[0]), .A2(sel[3]), .ZN(n80) );
  BUF_X1 U4 ( .A(n99), .Z(n101) );
  BUF_X1 U5 ( .A(n99), .Z(n100) );
  BUF_X1 U6 ( .A(n99), .Z(n102) );
  BUF_X1 U7 ( .A(n12), .Z(n88) );
  BUF_X1 U8 ( .A(n7), .Z(n103) );
  BUF_X1 U9 ( .A(n10), .Z(n93) );
  BUF_X1 U10 ( .A(n7), .Z(n104) );
  BUF_X1 U11 ( .A(n10), .Z(n94) );
  BUF_X1 U12 ( .A(n9), .Z(n98) );
  BUF_X1 U13 ( .A(n11), .Z(n92) );
  BUF_X1 U14 ( .A(n11), .Z(n90) );
  BUF_X1 U15 ( .A(n11), .Z(n91) );
  BUF_X1 U16 ( .A(n9), .Z(n96) );
  BUF_X1 U17 ( .A(n12), .Z(n87) );
  BUF_X1 U18 ( .A(n9), .Z(n97) );
  BUF_X1 U19 ( .A(n12), .Z(n89) );
  BUF_X1 U20 ( .A(n7), .Z(n105) );
  BUF_X1 U21 ( .A(n10), .Z(n95) );
  INV_X1 U22 ( .A(n83), .ZN(n78) );
  BUF_X1 U23 ( .A(n8), .Z(n99) );
  NOR4_X1 U24 ( .A1(n93), .A2(n96), .A3(n90), .A4(n83), .ZN(n8) );
  NAND2_X1 U25 ( .A1(n21), .A2(n22), .ZN(o[4]) );
  AOI222_X1 U26 ( .A1(out_sub[4]), .A2(n95), .B1(out_sr[4]), .B2(n90), .C1(
        out_cmp[4]), .C2(n87), .ZN(n21) );
  AOI222_X1 U27 ( .A1(out_sl[4]), .A2(n103), .B1(out_log[4]), .B2(n100), .C1(
        out_add[4]), .C2(n98), .ZN(n22) );
  NAND2_X1 U28 ( .A1(n5), .A2(n6), .ZN(o[9]) );
  AOI222_X1 U29 ( .A1(out_sub[9]), .A2(n95), .B1(out_sr[9]), .B2(n91), .C1(
        out_cmp[9]), .C2(n88), .ZN(n5) );
  AOI222_X1 U30 ( .A1(out_sl[9]), .A2(n104), .B1(out_log[9]), .B2(n100), .C1(
        out_add[9]), .C2(n98), .ZN(n6) );
  NAND2_X1 U31 ( .A1(n51), .A2(n52), .ZN(o[1]) );
  AOI222_X1 U32 ( .A1(out_sub[1]), .A2(n93), .B1(out_sr[1]), .B2(n91), .C1(
        out_cmp[1]), .C2(n88), .ZN(n51) );
  AOI222_X1 U33 ( .A1(out_sl[1]), .A2(n104), .B1(out_log[1]), .B2(n101), .C1(
        out_add[1]), .C2(n97), .ZN(n52) );
  NAND2_X1 U34 ( .A1(n29), .A2(n30), .ZN(o[2]) );
  AOI222_X1 U35 ( .A1(out_sub[2]), .A2(n94), .B1(out_sr[2]), .B2(n90), .C1(
        out_cmp[2]), .C2(n87), .ZN(n29) );
  AOI222_X1 U36 ( .A1(out_sl[2]), .A2(n103), .B1(out_log[2]), .B2(n100), .C1(
        out_add[2]), .C2(n97), .ZN(n30) );
  NAND2_X1 U37 ( .A1(n41), .A2(n42), .ZN(o[24]) );
  AOI222_X1 U38 ( .A1(out_sub[24]), .A2(n94), .B1(out_sr[24]), .B2(n91), .C1(
        out_cmp[24]), .C2(n88), .ZN(n41) );
  AOI222_X1 U39 ( .A1(out_sl[24]), .A2(n104), .B1(out_log[24]), .B2(n101), 
        .C1(out_add[24]), .C2(n97), .ZN(n42) );
  NOR2_X1 U40 ( .A1(n103), .A2(n76), .ZN(n75) );
  AOI221_X1 U41 ( .B1(out_sr[0]), .B2(n92), .C1(out_cmp[0]), .C2(n87), .A(n77), 
        .ZN(n76) );
  NOR3_X1 U42 ( .A1(n78), .A2(n87), .A3(n79), .ZN(n77) );
  AOI22_X1 U43 ( .A1(n80), .A2(n81), .B1(out_eq[0]), .B2(sel[3]), .ZN(n79) );
  NAND2_X1 U44 ( .A1(n71), .A2(n72), .ZN(o[10]) );
  AOI222_X1 U45 ( .A1(out_sub[10]), .A2(n93), .B1(out_sr[10]), .B2(n92), .C1(
        out_cmp[10]), .C2(n87), .ZN(n71) );
  AOI222_X1 U46 ( .A1(out_sl[10]), .A2(n103), .B1(out_log[10]), .B2(n102), 
        .C1(out_add[10]), .C2(n96), .ZN(n72) );
  NAND2_X1 U47 ( .A1(n69), .A2(n70), .ZN(o[11]) );
  AOI222_X1 U48 ( .A1(out_sub[11]), .A2(n93), .B1(out_sr[11]), .B2(n92), .C1(
        out_cmp[11]), .C2(n89), .ZN(n69) );
  AOI222_X1 U49 ( .A1(out_sl[11]), .A2(n105), .B1(out_log[11]), .B2(n102), 
        .C1(out_add[11]), .C2(n96), .ZN(n70) );
  NAND2_X1 U50 ( .A1(n67), .A2(n68), .ZN(o[12]) );
  AOI222_X1 U51 ( .A1(out_sub[12]), .A2(n93), .B1(out_sr[12]), .B2(n92), .C1(
        out_cmp[12]), .C2(n89), .ZN(n67) );
  AOI222_X1 U52 ( .A1(out_sl[12]), .A2(n105), .B1(out_log[12]), .B2(n102), 
        .C1(out_add[12]), .C2(n96), .ZN(n68) );
  NAND2_X1 U53 ( .A1(n65), .A2(n66), .ZN(o[13]) );
  AOI222_X1 U54 ( .A1(out_sub[13]), .A2(n93), .B1(out_sr[13]), .B2(n92), .C1(
        out_cmp[13]), .C2(n89), .ZN(n65) );
  AOI222_X1 U55 ( .A1(out_sl[13]), .A2(n105), .B1(out_log[13]), .B2(n102), 
        .C1(out_add[13]), .C2(n96), .ZN(n66) );
  NAND2_X1 U56 ( .A1(n63), .A2(n64), .ZN(o[14]) );
  AOI222_X1 U57 ( .A1(out_sub[14]), .A2(n93), .B1(out_sr[14]), .B2(n92), .C1(
        out_cmp[14]), .C2(n89), .ZN(n63) );
  AOI222_X1 U58 ( .A1(out_sl[14]), .A2(n105), .B1(out_log[14]), .B2(n102), 
        .C1(out_add[14]), .C2(n96), .ZN(n64) );
  NAND2_X1 U59 ( .A1(n61), .A2(n62), .ZN(o[15]) );
  AOI222_X1 U60 ( .A1(out_sub[15]), .A2(n93), .B1(out_sr[15]), .B2(n92), .C1(
        out_cmp[15]), .C2(n89), .ZN(n61) );
  AOI222_X1 U61 ( .A1(out_sl[15]), .A2(n105), .B1(out_log[15]), .B2(n102), 
        .C1(out_add[15]), .C2(n96), .ZN(n62) );
  NAND2_X1 U62 ( .A1(n59), .A2(n60), .ZN(o[16]) );
  AOI222_X1 U63 ( .A1(out_sub[16]), .A2(n93), .B1(out_sr[16]), .B2(n92), .C1(
        out_cmp[16]), .C2(n89), .ZN(n59) );
  AOI222_X1 U64 ( .A1(out_sl[16]), .A2(n105), .B1(out_log[16]), .B2(n102), 
        .C1(out_add[16]), .C2(n96), .ZN(n60) );
  NAND2_X1 U65 ( .A1(n57), .A2(n58), .ZN(o[17]) );
  AOI222_X1 U66 ( .A1(out_sub[17]), .A2(n93), .B1(out_sr[17]), .B2(n92), .C1(
        out_cmp[17]), .C2(n89), .ZN(n57) );
  AOI222_X1 U67 ( .A1(out_sl[17]), .A2(n105), .B1(out_log[17]), .B2(n101), 
        .C1(out_add[17]), .C2(n96), .ZN(n58) );
  NAND2_X1 U68 ( .A1(n23), .A2(n24), .ZN(o[3]) );
  AOI222_X1 U69 ( .A1(out_sub[3]), .A2(n95), .B1(out_sr[3]), .B2(n90), .C1(
        out_cmp[3]), .C2(n87), .ZN(n23) );
  AOI222_X1 U70 ( .A1(out_sl[3]), .A2(n103), .B1(out_log[3]), .B2(n100), .C1(
        out_add[3]), .C2(n98), .ZN(n24) );
  NAND2_X1 U71 ( .A1(n19), .A2(n20), .ZN(o[5]) );
  AOI222_X1 U72 ( .A1(out_sub[5]), .A2(n95), .B1(out_sr[5]), .B2(n90), .C1(
        out_cmp[5]), .C2(n87), .ZN(n19) );
  AOI222_X1 U73 ( .A1(out_sl[5]), .A2(n103), .B1(out_log[5]), .B2(n100), .C1(
        out_add[5]), .C2(n98), .ZN(n20) );
  NAND2_X1 U74 ( .A1(n17), .A2(n18), .ZN(o[6]) );
  AOI222_X1 U75 ( .A1(out_sub[6]), .A2(n95), .B1(out_sr[6]), .B2(n90), .C1(
        out_cmp[6]), .C2(n87), .ZN(n17) );
  AOI222_X1 U76 ( .A1(out_sl[6]), .A2(n103), .B1(out_log[6]), .B2(n100), .C1(
        out_add[6]), .C2(n98), .ZN(n18) );
  NAND2_X1 U77 ( .A1(n15), .A2(n16), .ZN(o[7]) );
  AOI222_X1 U78 ( .A1(out_sub[7]), .A2(n95), .B1(out_sr[7]), .B2(n90), .C1(
        out_cmp[7]), .C2(n87), .ZN(n15) );
  AOI222_X1 U79 ( .A1(out_sl[7]), .A2(n103), .B1(out_log[7]), .B2(n100), .C1(
        out_add[7]), .C2(n98), .ZN(n16) );
  NAND2_X1 U80 ( .A1(n13), .A2(n14), .ZN(o[8]) );
  AOI222_X1 U81 ( .A1(out_sub[8]), .A2(n95), .B1(out_sr[8]), .B2(n90), .C1(
        out_cmp[8]), .C2(n87), .ZN(n13) );
  AOI222_X1 U82 ( .A1(out_sl[8]), .A2(n103), .B1(out_log[8]), .B2(n100), .C1(
        out_add[8]), .C2(n98), .ZN(n14) );
  NAND2_X1 U83 ( .A1(n55), .A2(n56), .ZN(o[18]) );
  AOI222_X1 U84 ( .A1(out_sub[18]), .A2(n93), .B1(out_sr[18]), .B2(n91), .C1(
        out_cmp[18]), .C2(n89), .ZN(n55) );
  AOI222_X1 U85 ( .A1(out_sl[18]), .A2(n104), .B1(out_log[18]), .B2(n101), 
        .C1(out_add[18]), .C2(n96), .ZN(n56) );
  NAND2_X1 U86 ( .A1(n53), .A2(n54), .ZN(o[19]) );
  AOI222_X1 U87 ( .A1(out_sub[19]), .A2(n93), .B1(out_sr[19]), .B2(n91), .C1(
        out_cmp[19]), .C2(n88), .ZN(n53) );
  AOI222_X1 U88 ( .A1(out_sl[19]), .A2(n104), .B1(out_log[19]), .B2(n101), 
        .C1(out_add[19]), .C2(n96), .ZN(n54) );
  NAND2_X1 U89 ( .A1(n49), .A2(n50), .ZN(o[20]) );
  AOI222_X1 U90 ( .A1(out_sub[20]), .A2(n94), .B1(out_sr[20]), .B2(n91), .C1(
        out_cmp[20]), .C2(n88), .ZN(n49) );
  AOI222_X1 U91 ( .A1(out_sl[20]), .A2(n104), .B1(out_log[20]), .B2(n101), 
        .C1(out_add[20]), .C2(n97), .ZN(n50) );
  NAND2_X1 U92 ( .A1(n47), .A2(n48), .ZN(o[21]) );
  AOI222_X1 U93 ( .A1(out_sub[21]), .A2(n94), .B1(out_sr[21]), .B2(n91), .C1(
        out_cmp[21]), .C2(n88), .ZN(n47) );
  AOI222_X1 U94 ( .A1(out_sl[21]), .A2(n104), .B1(out_log[21]), .B2(n101), 
        .C1(out_add[21]), .C2(n97), .ZN(n48) );
  NAND2_X1 U95 ( .A1(n45), .A2(n46), .ZN(o[22]) );
  AOI222_X1 U96 ( .A1(out_sub[22]), .A2(n94), .B1(out_sr[22]), .B2(n91), .C1(
        out_cmp[22]), .C2(n88), .ZN(n45) );
  AOI222_X1 U97 ( .A1(out_sl[22]), .A2(n104), .B1(out_log[22]), .B2(n101), 
        .C1(out_add[22]), .C2(n97), .ZN(n46) );
  NAND2_X1 U98 ( .A1(n43), .A2(n44), .ZN(o[23]) );
  AOI222_X1 U99 ( .A1(out_sub[23]), .A2(n94), .B1(out_sr[23]), .B2(n91), .C1(
        out_cmp[23]), .C2(n88), .ZN(n43) );
  AOI222_X1 U100 ( .A1(out_sl[23]), .A2(n104), .B1(out_log[23]), .B2(n101), 
        .C1(out_add[23]), .C2(n97), .ZN(n44) );
  NAND2_X1 U101 ( .A1(n39), .A2(n40), .ZN(o[25]) );
  AOI222_X1 U102 ( .A1(out_sub[25]), .A2(n94), .B1(out_sr[25]), .B2(n91), .C1(
        out_cmp[25]), .C2(n88), .ZN(n39) );
  AOI222_X1 U103 ( .A1(out_sl[25]), .A2(n104), .B1(out_log[25]), .B2(n101), 
        .C1(out_add[25]), .C2(n97), .ZN(n40) );
  NAND2_X1 U104 ( .A1(n37), .A2(n38), .ZN(o[26]) );
  AOI222_X1 U105 ( .A1(out_sub[26]), .A2(n94), .B1(out_sr[26]), .B2(n91), .C1(
        out_cmp[26]), .C2(n88), .ZN(n37) );
  AOI222_X1 U106 ( .A1(out_sl[26]), .A2(n104), .B1(out_log[26]), .B2(n101), 
        .C1(out_add[26]), .C2(n97), .ZN(n38) );
  NAND2_X1 U107 ( .A1(n35), .A2(n36), .ZN(o[27]) );
  AOI222_X1 U108 ( .A1(out_sub[27]), .A2(n94), .B1(out_sr[27]), .B2(n91), .C1(
        out_cmp[27]), .C2(n88), .ZN(n35) );
  AOI222_X1 U109 ( .A1(out_sl[27]), .A2(n104), .B1(out_log[27]), .B2(n101), 
        .C1(out_add[27]), .C2(n97), .ZN(n36) );
  NAND2_X1 U110 ( .A1(n33), .A2(n34), .ZN(o[28]) );
  AOI222_X1 U111 ( .A1(out_sub[28]), .A2(n94), .B1(out_sr[28]), .B2(n90), .C1(
        out_cmp[28]), .C2(n88), .ZN(n33) );
  AOI222_X1 U112 ( .A1(out_sl[28]), .A2(n104), .B1(out_log[28]), .B2(n100), 
        .C1(out_add[28]), .C2(n97), .ZN(n34) );
  NAND2_X1 U113 ( .A1(n31), .A2(n32), .ZN(o[29]) );
  AOI222_X1 U114 ( .A1(out_sub[29]), .A2(n94), .B1(out_sr[29]), .B2(n90), .C1(
        out_cmp[29]), .C2(n88), .ZN(n31) );
  AOI222_X1 U115 ( .A1(out_sl[29]), .A2(n103), .B1(out_log[29]), .B2(n100), 
        .C1(out_add[29]), .C2(n97), .ZN(n32) );
  NAND2_X1 U116 ( .A1(n27), .A2(n28), .ZN(o[30]) );
  AOI222_X1 U117 ( .A1(out_sub[30]), .A2(n94), .B1(out_sr[30]), .B2(n90), .C1(
        out_cmp[30]), .C2(n87), .ZN(n27) );
  AOI222_X1 U118 ( .A1(out_sl[30]), .A2(n103), .B1(out_log[30]), .B2(n100), 
        .C1(out_add[30]), .C2(n98), .ZN(n28) );
  NAND2_X1 U119 ( .A1(n25), .A2(n26), .ZN(o[31]) );
  AOI222_X1 U120 ( .A1(out_sub[31]), .A2(n94), .B1(out_sr[31]), .B2(n90), .C1(
        out_cmp[31]), .C2(n87), .ZN(n25) );
  AOI222_X1 U121 ( .A1(out_sl[31]), .A2(n103), .B1(out_log[31]), .B2(n100), 
        .C1(out_add[31]), .C2(n98), .ZN(n26) );
  NAND2_X1 U122 ( .A1(n73), .A2(n74), .ZN(o[0]) );
  AOI22_X1 U123 ( .A1(out_add[0]), .A2(n96), .B1(out_sub[0]), .B2(n93), .ZN(
        n73) );
  AOI221_X1 U124 ( .B1(out_log[0]), .B2(n102), .C1(out_sl[0]), .C2(n103), .A(
        n75), .ZN(n74) );
  NOR4_X1 U125 ( .A1(sel[0]), .A2(sel[1]), .A3(sel[2]), .A4(sel[3]), .ZN(n9)
         );
  NOR3_X1 U126 ( .A1(sel[0]), .A2(sel[3]), .A3(n78), .ZN(n7) );
  NOR3_X1 U127 ( .A1(n107), .A2(sel[0]), .A3(n78), .ZN(n12) );
  NOR2_X1 U128 ( .A1(n106), .A2(sel[2]), .ZN(n83) );
  AND3_X1 U129 ( .A1(n106), .A2(n107), .A3(sel[2]), .ZN(n11) );
  AND4_X1 U130 ( .A1(sel[3]), .A2(sel[0]), .A3(sel[2]), .A4(sel[1]), .ZN(n10)
         );
  INV_X1 U131 ( .A(sel[1]), .ZN(n106) );
  INV_X1 U132 ( .A(sel[3]), .ZN(n107) );
endmodule


module logic_n_n32 ( r1, r2, s0, s1, s2, s3, y );
  input [31:0] r1;
  input [31:0] r2;
  output [31:0] y;
  input s0, s1, s2, s3;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  logic_0 logic_i_0 ( .r1(r1[0]), .r2(r2[0]), .s0(n3), .s1(n6), .s2(n9), .s3(
        n12), .y(y[0]) );
  logic_31 logic_i_1 ( .r1(r1[1]), .r2(r2[1]), .s0(n1), .s1(n4), .s2(n7), .s3(
        n10), .y(y[1]) );
  logic_30 logic_i_2 ( .r1(r1[2]), .r2(r2[2]), .s0(n1), .s1(n4), .s2(n7), .s3(
        n10), .y(y[2]) );
  logic_29 logic_i_3 ( .r1(r1[3]), .r2(r2[3]), .s0(n1), .s1(n4), .s2(n7), .s3(
        n10), .y(y[3]) );
  logic_28 logic_i_4 ( .r1(r1[4]), .r2(r2[4]), .s0(n1), .s1(n4), .s2(n7), .s3(
        n10), .y(y[4]) );
  logic_27 logic_i_5 ( .r1(r1[5]), .r2(r2[5]), .s0(n1), .s1(n4), .s2(n7), .s3(
        n10), .y(y[5]) );
  logic_26 logic_i_6 ( .r1(r1[6]), .r2(r2[6]), .s0(n1), .s1(n4), .s2(n7), .s3(
        n10), .y(y[6]) );
  logic_25 logic_i_7 ( .r1(r1[7]), .r2(r2[7]), .s0(n1), .s1(n4), .s2(n7), .s3(
        n10), .y(y[7]) );
  logic_24 logic_i_8 ( .r1(r1[8]), .r2(r2[8]), .s0(n1), .s1(n4), .s2(n7), .s3(
        n10), .y(y[8]) );
  logic_23 logic_i_9 ( .r1(r1[9]), .r2(r2[9]), .s0(n1), .s1(n4), .s2(n7), .s3(
        n10), .y(y[9]) );
  logic_22 logic_i_10 ( .r1(r1[10]), .r2(r2[10]), .s0(n1), .s1(n4), .s2(n7), 
        .s3(n10), .y(y[10]) );
  logic_21 logic_i_11 ( .r1(r1[11]), .r2(r2[11]), .s0(n1), .s1(n4), .s2(n7), 
        .s3(n10), .y(y[11]) );
  logic_20 logic_i_12 ( .r1(r1[12]), .r2(r2[12]), .s0(n1), .s1(n4), .s2(n7), 
        .s3(n10), .y(y[12]) );
  logic_19 logic_i_13 ( .r1(r1[13]), .r2(r2[13]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[13]) );
  logic_18 logic_i_14 ( .r1(r1[14]), .r2(r2[14]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[14]) );
  logic_17 logic_i_15 ( .r1(r1[15]), .r2(r2[15]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[15]) );
  logic_16 logic_i_16 ( .r1(r1[16]), .r2(r2[16]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[16]) );
  logic_15 logic_i_17 ( .r1(r1[17]), .r2(r2[17]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[17]) );
  logic_14 logic_i_18 ( .r1(r1[18]), .r2(r2[18]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[18]) );
  logic_13 logic_i_19 ( .r1(r1[19]), .r2(r2[19]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[19]) );
  logic_12 logic_i_20 ( .r1(r1[20]), .r2(r2[20]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[20]) );
  logic_11 logic_i_21 ( .r1(r1[21]), .r2(r2[21]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[21]) );
  logic_10 logic_i_22 ( .r1(r1[22]), .r2(r2[22]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[22]) );
  logic_9 logic_i_23 ( .r1(r1[23]), .r2(r2[23]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[23]) );
  logic_8 logic_i_24 ( .r1(r1[24]), .r2(r2[24]), .s0(n2), .s1(n5), .s2(n8), 
        .s3(n11), .y(y[24]) );
  logic_7 logic_i_25 ( .r1(r1[25]), .r2(r2[25]), .s0(n3), .s1(n6), .s2(n9), 
        .s3(n12), .y(y[25]) );
  logic_6 logic_i_26 ( .r1(r1[26]), .r2(r2[26]), .s0(n3), .s1(n6), .s2(n9), 
        .s3(n12), .y(y[26]) );
  logic_5 logic_i_27 ( .r1(r1[27]), .r2(r2[27]), .s0(n3), .s1(n6), .s2(n9), 
        .s3(n12), .y(y[27]) );
  logic_4 logic_i_28 ( .r1(r1[28]), .r2(r2[28]), .s0(n3), .s1(n6), .s2(n9), 
        .s3(n12), .y(y[28]) );
  logic_3 logic_i_29 ( .r1(r1[29]), .r2(r2[29]), .s0(n3), .s1(n6), .s2(n9), 
        .s3(n12), .y(y[29]) );
  logic_2 logic_i_30 ( .r1(r1[30]), .r2(r2[30]), .s0(n3), .s1(n6), .s2(n9), 
        .s3(n12), .y(y[30]) );
  logic_1 logic_i_31 ( .r1(r1[31]), .r2(r2[31]), .s0(n3), .s1(n6), .s2(n9), 
        .s3(n12), .y(y[31]) );
  BUF_X1 U1 ( .A(s0), .Z(n1) );
  BUF_X1 U2 ( .A(s0), .Z(n2) );
  BUF_X1 U3 ( .A(s2), .Z(n7) );
  BUF_X1 U4 ( .A(s2), .Z(n8) );
  BUF_X1 U5 ( .A(s1), .Z(n4) );
  BUF_X1 U6 ( .A(s1), .Z(n5) );
  BUF_X1 U7 ( .A(s3), .Z(n10) );
  BUF_X1 U8 ( .A(s3), .Z(n11) );
  BUF_X1 U9 ( .A(s0), .Z(n3) );
  BUF_X1 U10 ( .A(s1), .Z(n6) );
  BUF_X1 U11 ( .A(s2), .Z(n9) );
  BUF_X1 U12 ( .A(s3), .Z(n12) );
endmodule


module xor_2_353 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module comparator_n32 ( a, b, cout, z );
  input [31:0] a;
  input [31:0] b;
  output cout, z;

  wire   [31:0] b_not;
  wire   [31:0] s;

  not_n_n32_1 b_negate ( .a(b), .y(b_not) );
  rca_n_n32_1 sub ( .a(a), .b(b_not), .c_in(1'b1), .sum(s), .c_out(cout) );
  nor_n1_n32 big_nor ( .a(s), .y(z) );
endmodule


module barrel_shifter_right_n32 ( x, pos, shift_type, y );
  input [31:0] x;
  input [4:0] pos;
  output [31:0] y;
  input shift_type;
  wire   \temp[4][31] , \temp[4][30] , \temp[4][29] , \temp[4][28] ,
         \temp[4][27] , \temp[4][26] , \temp[4][25] , \temp[4][24] ,
         \temp[4][23] , \temp[4][22] , \temp[4][21] , \temp[4][20] ,
         \temp[4][19] , \temp[4][18] , \temp[4][17] , \temp[4][16] ,
         \temp[4][15] , \temp[4][14] , \temp[4][13] , \temp[4][12] ,
         \temp[4][11] , \temp[4][10] , \temp[4][9] , \temp[4][8] ,
         \temp[4][7] , \temp[4][6] , \temp[4][5] , \temp[4][4] , \temp[4][3] ,
         \temp[4][2] , \temp[4][1] , \temp[4][0] , \temp[3][31] ,
         \temp[3][30] , \temp[3][29] , \temp[3][28] , \temp[3][27] ,
         \temp[3][26] , \temp[3][25] , \temp[3][24] , \temp[3][23] ,
         \temp[3][22] , \temp[3][21] , \temp[3][20] , \temp[3][19] ,
         \temp[3][18] , \temp[3][17] , \temp[3][16] , \temp[3][15] ,
         \temp[3][14] , \temp[3][13] , \temp[3][12] , \temp[3][11] ,
         \temp[3][10] , \temp[3][9] , \temp[3][8] , \temp[3][7] , \temp[3][6] ,
         \temp[3][5] , \temp[3][4] , \temp[3][3] , \temp[3][2] , \temp[3][1] ,
         \temp[3][0] , \temp[2][31] , \temp[2][30] , \temp[2][29] ,
         \temp[2][28] , \temp[2][27] , \temp[2][26] , \temp[2][25] ,
         \temp[2][24] , \temp[2][23] , \temp[2][22] , \temp[2][21] ,
         \temp[2][20] , \temp[2][19] , \temp[2][18] , \temp[2][17] ,
         \temp[2][16] , \temp[2][15] , \temp[2][14] , \temp[2][13] ,
         \temp[2][12] , \temp[2][11] , \temp[2][10] , \temp[2][9] ,
         \temp[2][8] , \temp[2][7] , \temp[2][6] , \temp[2][5] , \temp[2][4] ,
         \temp[2][3] , \temp[2][2] , \temp[2][1] , \temp[2][0] , \temp[1][31] ,
         \temp[1][30] , \temp[1][29] , \temp[1][28] , \temp[1][27] ,
         \temp[1][26] , \temp[1][25] , \temp[1][24] , \temp[1][23] ,
         \temp[1][22] , \temp[1][21] , \temp[1][20] , \temp[1][19] ,
         \temp[1][18] , \temp[1][17] , \temp[1][16] , \temp[1][15] ,
         \temp[1][14] , \temp[1][13] , \temp[1][12] , \temp[1][11] ,
         \temp[1][10] , \temp[1][9] , \temp[1][8] , \temp[1][7] , \temp[1][6] ,
         \temp[1][5] , \temp[1][4] , \temp[1][3] , \temp[1][2] , \temp[1][1] ,
         \temp[1][0] , n3, n6, n9, n12, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33;
  tri   [31:0] y;
  assign n3 = pos[0];
  assign n6 = pos[1];
  assign n9 = pos[2];
  assign n12 = pos[3];
  assign n15 = pos[4];

  mux21_192 mux21_k_0_0 ( .a(x[0]), .b(x[1]), .s(n19), .y(\temp[1][0] ) );
  mux21_191 mux21_k_0_1 ( .a(x[1]), .b(x[2]), .s(n19), .y(\temp[1][1] ) );
  mux21_190 mux21_k_0_2 ( .a(x[2]), .b(x[3]), .s(n19), .y(\temp[1][2] ) );
  mux21_189 mux21_k_0_3 ( .a(x[3]), .b(x[4]), .s(n19), .y(\temp[1][3] ) );
  mux21_188 mux21_k_0_4 ( .a(x[4]), .b(x[5]), .s(n19), .y(\temp[1][4] ) );
  mux21_187 mux21_k_0_5 ( .a(x[5]), .b(x[6]), .s(n19), .y(\temp[1][5] ) );
  mux21_186 mux21_k_0_6 ( .a(x[6]), .b(x[7]), .s(n19), .y(\temp[1][6] ) );
  mux21_185 mux21_k_0_7 ( .a(x[7]), .b(x[8]), .s(n19), .y(\temp[1][7] ) );
  mux21_184 mux21_k_0_8 ( .a(x[8]), .b(x[9]), .s(n19), .y(\temp[1][8] ) );
  mux21_183 mux21_k_0_9 ( .a(x[9]), .b(x[10]), .s(n19), .y(\temp[1][9] ) );
  mux21_182 mux21_k_0_10 ( .a(x[10]), .b(x[11]), .s(n19), .y(\temp[1][10] ) );
  mux21_181 mux21_k_0_11 ( .a(x[11]), .b(x[12]), .s(n19), .y(\temp[1][11] ) );
  mux21_180 mux21_k_0_12 ( .a(x[12]), .b(x[13]), .s(n20), .y(\temp[1][12] ) );
  mux21_179 mux21_k_0_13 ( .a(x[13]), .b(x[14]), .s(n20), .y(\temp[1][13] ) );
  mux21_178 mux21_k_0_14 ( .a(x[14]), .b(x[15]), .s(n20), .y(\temp[1][14] ) );
  mux21_177 mux21_k_0_15 ( .a(x[15]), .b(x[16]), .s(n20), .y(\temp[1][15] ) );
  mux21_176 mux21_k_0_16 ( .a(x[16]), .b(x[17]), .s(n20), .y(\temp[1][16] ) );
  mux21_175 mux21_k_0_17 ( .a(x[17]), .b(x[18]), .s(n20), .y(\temp[1][17] ) );
  mux21_174 mux21_k_0_18 ( .a(x[18]), .b(x[19]), .s(n20), .y(\temp[1][18] ) );
  mux21_173 mux21_k_0_19 ( .a(x[19]), .b(x[20]), .s(n20), .y(\temp[1][19] ) );
  mux21_172 mux21_k_0_20 ( .a(x[20]), .b(x[21]), .s(n20), .y(\temp[1][20] ) );
  mux21_171 mux21_k_0_21 ( .a(x[21]), .b(x[22]), .s(n20), .y(\temp[1][21] ) );
  mux21_170 mux21_k_0_22 ( .a(x[22]), .b(x[23]), .s(n20), .y(\temp[1][22] ) );
  mux21_169 mux21_k_0_23 ( .a(x[23]), .b(x[24]), .s(n20), .y(\temp[1][23] ) );
  mux21_168 mux21_k_0_24 ( .a(x[24]), .b(x[25]), .s(n21), .y(\temp[1][24] ) );
  mux21_167 mux21_k_0_25 ( .a(x[25]), .b(x[26]), .s(n21), .y(\temp[1][25] ) );
  mux21_166 mux21_k_0_26 ( .a(x[26]), .b(x[27]), .s(n21), .y(\temp[1][26] ) );
  mux21_165 mux21_k_0_27 ( .a(x[27]), .b(x[28]), .s(n21), .y(\temp[1][27] ) );
  mux21_164 mux21_k_0_28 ( .a(x[28]), .b(x[29]), .s(n21), .y(\temp[1][28] ) );
  mux21_163 mux21_k_0_29 ( .a(x[29]), .b(x[30]), .s(n21), .y(\temp[1][29] ) );
  mux21_162 mux21_k_0_30 ( .a(x[30]), .b(x[31]), .s(n21), .y(\temp[1][30] ) );
  mux21_161 mux21_j_0_0 ( .a(x[31]), .b(n16), .s(n21), .y(\temp[1][31] ) );
  mux21_160 mux21_k_1_0 ( .a(\temp[1][0] ), .b(\temp[1][2] ), .s(n22), .y(
        \temp[2][0] ) );
  mux21_159 mux21_k_1_1 ( .a(\temp[1][1] ), .b(\temp[1][3] ), .s(n22), .y(
        \temp[2][1] ) );
  mux21_158 mux21_k_1_2 ( .a(\temp[1][2] ), .b(\temp[1][4] ), .s(n22), .y(
        \temp[2][2] ) );
  mux21_157 mux21_k_1_3 ( .a(\temp[1][3] ), .b(\temp[1][5] ), .s(n22), .y(
        \temp[2][3] ) );
  mux21_156 mux21_k_1_4 ( .a(\temp[1][4] ), .b(\temp[1][6] ), .s(n22), .y(
        \temp[2][4] ) );
  mux21_155 mux21_k_1_5 ( .a(\temp[1][5] ), .b(\temp[1][7] ), .s(n22), .y(
        \temp[2][5] ) );
  mux21_154 mux21_k_1_6 ( .a(\temp[1][6] ), .b(\temp[1][8] ), .s(n22), .y(
        \temp[2][6] ) );
  mux21_153 mux21_k_1_7 ( .a(\temp[1][7] ), .b(\temp[1][9] ), .s(n22), .y(
        \temp[2][7] ) );
  mux21_152 mux21_k_1_8 ( .a(\temp[1][8] ), .b(\temp[1][10] ), .s(n22), .y(
        \temp[2][8] ) );
  mux21_151 mux21_k_1_9 ( .a(\temp[1][9] ), .b(\temp[1][11] ), .s(n22), .y(
        \temp[2][9] ) );
  mux21_150 mux21_k_1_10 ( .a(\temp[1][10] ), .b(\temp[1][12] ), .s(n22), .y(
        \temp[2][10] ) );
  mux21_149 mux21_k_1_11 ( .a(\temp[1][11] ), .b(\temp[1][13] ), .s(n22), .y(
        \temp[2][11] ) );
  mux21_148 mux21_k_1_12 ( .a(\temp[1][12] ), .b(\temp[1][14] ), .s(n23), .y(
        \temp[2][12] ) );
  mux21_147 mux21_k_1_13 ( .a(\temp[1][13] ), .b(\temp[1][15] ), .s(n23), .y(
        \temp[2][13] ) );
  mux21_146 mux21_k_1_14 ( .a(\temp[1][14] ), .b(\temp[1][16] ), .s(n23), .y(
        \temp[2][14] ) );
  mux21_145 mux21_k_1_15 ( .a(\temp[1][15] ), .b(\temp[1][17] ), .s(n23), .y(
        \temp[2][15] ) );
  mux21_144 mux21_k_1_16 ( .a(\temp[1][16] ), .b(\temp[1][18] ), .s(n23), .y(
        \temp[2][16] ) );
  mux21_143 mux21_k_1_17 ( .a(\temp[1][17] ), .b(\temp[1][19] ), .s(n23), .y(
        \temp[2][17] ) );
  mux21_142 mux21_k_1_18 ( .a(\temp[1][18] ), .b(\temp[1][20] ), .s(n23), .y(
        \temp[2][18] ) );
  mux21_141 mux21_k_1_19 ( .a(\temp[1][19] ), .b(\temp[1][21] ), .s(n23), .y(
        \temp[2][19] ) );
  mux21_140 mux21_k_1_20 ( .a(\temp[1][20] ), .b(\temp[1][22] ), .s(n23), .y(
        \temp[2][20] ) );
  mux21_139 mux21_k_1_21 ( .a(\temp[1][21] ), .b(\temp[1][23] ), .s(n23), .y(
        \temp[2][21] ) );
  mux21_138 mux21_k_1_22 ( .a(\temp[1][22] ), .b(\temp[1][24] ), .s(n23), .y(
        \temp[2][22] ) );
  mux21_137 mux21_k_1_23 ( .a(\temp[1][23] ), .b(\temp[1][25] ), .s(n23), .y(
        \temp[2][23] ) );
  mux21_136 mux21_k_1_24 ( .a(\temp[1][24] ), .b(\temp[1][26] ), .s(n24), .y(
        \temp[2][24] ) );
  mux21_135 mux21_k_1_25 ( .a(\temp[1][25] ), .b(\temp[1][27] ), .s(n24), .y(
        \temp[2][25] ) );
  mux21_134 mux21_k_1_26 ( .a(\temp[1][26] ), .b(\temp[1][28] ), .s(n24), .y(
        \temp[2][26] ) );
  mux21_133 mux21_k_1_27 ( .a(\temp[1][27] ), .b(\temp[1][29] ), .s(n24), .y(
        \temp[2][27] ) );
  mux21_132 mux21_k_1_28 ( .a(\temp[1][28] ), .b(\temp[1][30] ), .s(n24), .y(
        \temp[2][28] ) );
  mux21_131 mux21_k_1_29 ( .a(\temp[1][29] ), .b(\temp[1][31] ), .s(n24), .y(
        \temp[2][29] ) );
  mux21_130 mux21_j_1_0 ( .a(\temp[1][30] ), .b(n16), .s(n24), .y(
        \temp[2][30] ) );
  mux21_129 mux21_j_1_1 ( .a(\temp[1][31] ), .b(n16), .s(n24), .y(
        \temp[2][31] ) );
  mux21_128 mux21_k_2_0 ( .a(\temp[2][0] ), .b(\temp[2][4] ), .s(n25), .y(
        \temp[3][0] ) );
  mux21_127 mux21_k_2_1 ( .a(\temp[2][1] ), .b(\temp[2][5] ), .s(n25), .y(
        \temp[3][1] ) );
  mux21_126 mux21_k_2_2 ( .a(\temp[2][2] ), .b(\temp[2][6] ), .s(n25), .y(
        \temp[3][2] ) );
  mux21_125 mux21_k_2_3 ( .a(\temp[2][3] ), .b(\temp[2][7] ), .s(n25), .y(
        \temp[3][3] ) );
  mux21_124 mux21_k_2_4 ( .a(\temp[2][4] ), .b(\temp[2][8] ), .s(n25), .y(
        \temp[3][4] ) );
  mux21_123 mux21_k_2_5 ( .a(\temp[2][5] ), .b(\temp[2][9] ), .s(n25), .y(
        \temp[3][5] ) );
  mux21_122 mux21_k_2_6 ( .a(\temp[2][6] ), .b(\temp[2][10] ), .s(n25), .y(
        \temp[3][6] ) );
  mux21_121 mux21_k_2_7 ( .a(\temp[2][7] ), .b(\temp[2][11] ), .s(n25), .y(
        \temp[3][7] ) );
  mux21_120 mux21_k_2_8 ( .a(\temp[2][8] ), .b(\temp[2][12] ), .s(n25), .y(
        \temp[3][8] ) );
  mux21_119 mux21_k_2_9 ( .a(\temp[2][9] ), .b(\temp[2][13] ), .s(n25), .y(
        \temp[3][9] ) );
  mux21_118 mux21_k_2_10 ( .a(\temp[2][10] ), .b(\temp[2][14] ), .s(n25), .y(
        \temp[3][10] ) );
  mux21_117 mux21_k_2_11 ( .a(\temp[2][11] ), .b(\temp[2][15] ), .s(n25), .y(
        \temp[3][11] ) );
  mux21_116 mux21_k_2_12 ( .a(\temp[2][12] ), .b(\temp[2][16] ), .s(n26), .y(
        \temp[3][12] ) );
  mux21_115 mux21_k_2_13 ( .a(\temp[2][13] ), .b(\temp[2][17] ), .s(n26), .y(
        \temp[3][13] ) );
  mux21_114 mux21_k_2_14 ( .a(\temp[2][14] ), .b(\temp[2][18] ), .s(n26), .y(
        \temp[3][14] ) );
  mux21_113 mux21_k_2_15 ( .a(\temp[2][15] ), .b(\temp[2][19] ), .s(n26), .y(
        \temp[3][15] ) );
  mux21_112 mux21_k_2_16 ( .a(\temp[2][16] ), .b(\temp[2][20] ), .s(n26), .y(
        \temp[3][16] ) );
  mux21_111 mux21_k_2_17 ( .a(\temp[2][17] ), .b(\temp[2][21] ), .s(n26), .y(
        \temp[3][17] ) );
  mux21_110 mux21_k_2_18 ( .a(\temp[2][18] ), .b(\temp[2][22] ), .s(n26), .y(
        \temp[3][18] ) );
  mux21_109 mux21_k_2_19 ( .a(\temp[2][19] ), .b(\temp[2][23] ), .s(n26), .y(
        \temp[3][19] ) );
  mux21_108 mux21_k_2_20 ( .a(\temp[2][20] ), .b(\temp[2][24] ), .s(n26), .y(
        \temp[3][20] ) );
  mux21_107 mux21_k_2_21 ( .a(\temp[2][21] ), .b(\temp[2][25] ), .s(n26), .y(
        \temp[3][21] ) );
  mux21_106 mux21_k_2_22 ( .a(\temp[2][22] ), .b(\temp[2][26] ), .s(n26), .y(
        \temp[3][22] ) );
  mux21_105 mux21_k_2_23 ( .a(\temp[2][23] ), .b(\temp[2][27] ), .s(n26), .y(
        \temp[3][23] ) );
  mux21_104 mux21_k_2_24 ( .a(\temp[2][24] ), .b(\temp[2][28] ), .s(n27), .y(
        \temp[3][24] ) );
  mux21_103 mux21_k_2_25 ( .a(\temp[2][25] ), .b(\temp[2][29] ), .s(n27), .y(
        \temp[3][25] ) );
  mux21_102 mux21_k_2_26 ( .a(\temp[2][26] ), .b(\temp[2][30] ), .s(n27), .y(
        \temp[3][26] ) );
  mux21_101 mux21_k_2_27 ( .a(\temp[2][27] ), .b(\temp[2][31] ), .s(n27), .y(
        \temp[3][27] ) );
  mux21_100 mux21_j_2_0 ( .a(\temp[2][28] ), .b(n16), .s(n27), .y(
        \temp[3][28] ) );
  mux21_99 mux21_j_2_1 ( .a(\temp[2][29] ), .b(n16), .s(n27), .y(\temp[3][29] ) );
  mux21_98 mux21_j_2_2 ( .a(\temp[2][30] ), .b(n16), .s(n27), .y(\temp[3][30] ) );
  mux21_97 mux21_j_2_3 ( .a(\temp[2][31] ), .b(n16), .s(n27), .y(\temp[3][31] ) );
  mux21_96 mux21_k_3_0 ( .a(\temp[3][0] ), .b(\temp[3][8] ), .s(n28), .y(
        \temp[4][0] ) );
  mux21_95 mux21_k_3_1 ( .a(\temp[3][1] ), .b(\temp[3][9] ), .s(n28), .y(
        \temp[4][1] ) );
  mux21_94 mux21_k_3_2 ( .a(\temp[3][2] ), .b(\temp[3][10] ), .s(n28), .y(
        \temp[4][2] ) );
  mux21_93 mux21_k_3_3 ( .a(\temp[3][3] ), .b(\temp[3][11] ), .s(n28), .y(
        \temp[4][3] ) );
  mux21_92 mux21_k_3_4 ( .a(\temp[3][4] ), .b(\temp[3][12] ), .s(n28), .y(
        \temp[4][4] ) );
  mux21_91 mux21_k_3_5 ( .a(\temp[3][5] ), .b(\temp[3][13] ), .s(n28), .y(
        \temp[4][5] ) );
  mux21_90 mux21_k_3_6 ( .a(\temp[3][6] ), .b(\temp[3][14] ), .s(n28), .y(
        \temp[4][6] ) );
  mux21_89 mux21_k_3_7 ( .a(\temp[3][7] ), .b(\temp[3][15] ), .s(n28), .y(
        \temp[4][7] ) );
  mux21_88 mux21_k_3_8 ( .a(\temp[3][8] ), .b(\temp[3][16] ), .s(n28), .y(
        \temp[4][8] ) );
  mux21_87 mux21_k_3_9 ( .a(\temp[3][9] ), .b(\temp[3][17] ), .s(n28), .y(
        \temp[4][9] ) );
  mux21_86 mux21_k_3_10 ( .a(\temp[3][10] ), .b(\temp[3][18] ), .s(n28), .y(
        \temp[4][10] ) );
  mux21_85 mux21_k_3_11 ( .a(\temp[3][11] ), .b(\temp[3][19] ), .s(n28), .y(
        \temp[4][11] ) );
  mux21_84 mux21_k_3_12 ( .a(\temp[3][12] ), .b(\temp[3][20] ), .s(n29), .y(
        \temp[4][12] ) );
  mux21_83 mux21_k_3_13 ( .a(\temp[3][13] ), .b(\temp[3][21] ), .s(n29), .y(
        \temp[4][13] ) );
  mux21_82 mux21_k_3_14 ( .a(\temp[3][14] ), .b(\temp[3][22] ), .s(n29), .y(
        \temp[4][14] ) );
  mux21_81 mux21_k_3_15 ( .a(\temp[3][15] ), .b(\temp[3][23] ), .s(n29), .y(
        \temp[4][15] ) );
  mux21_80 mux21_k_3_16 ( .a(\temp[3][16] ), .b(\temp[3][24] ), .s(n29), .y(
        \temp[4][16] ) );
  mux21_79 mux21_k_3_17 ( .a(\temp[3][17] ), .b(\temp[3][25] ), .s(n29), .y(
        \temp[4][17] ) );
  mux21_78 mux21_k_3_18 ( .a(\temp[3][18] ), .b(\temp[3][26] ), .s(n29), .y(
        \temp[4][18] ) );
  mux21_77 mux21_k_3_19 ( .a(\temp[3][19] ), .b(\temp[3][27] ), .s(n29), .y(
        \temp[4][19] ) );
  mux21_76 mux21_k_3_20 ( .a(\temp[3][20] ), .b(\temp[3][28] ), .s(n29), .y(
        \temp[4][20] ) );
  mux21_75 mux21_k_3_21 ( .a(\temp[3][21] ), .b(\temp[3][29] ), .s(n29), .y(
        \temp[4][21] ) );
  mux21_74 mux21_k_3_22 ( .a(\temp[3][22] ), .b(\temp[3][30] ), .s(n29), .y(
        \temp[4][22] ) );
  mux21_73 mux21_k_3_23 ( .a(\temp[3][23] ), .b(\temp[3][31] ), .s(n29), .y(
        \temp[4][23] ) );
  mux21_72 mux21_j_3_0 ( .a(\temp[3][24] ), .b(n16), .s(n30), .y(\temp[4][24] ) );
  mux21_71 mux21_j_3_1 ( .a(\temp[3][25] ), .b(n16), .s(n30), .y(\temp[4][25] ) );
  mux21_70 mux21_j_3_2 ( .a(\temp[3][26] ), .b(n16), .s(n30), .y(\temp[4][26] ) );
  mux21_69 mux21_j_3_3 ( .a(\temp[3][27] ), .b(n16), .s(n30), .y(\temp[4][27] ) );
  mux21_68 mux21_j_3_4 ( .a(\temp[3][28] ), .b(n16), .s(n30), .y(\temp[4][28] ) );
  mux21_67 mux21_j_3_5 ( .a(\temp[3][29] ), .b(n17), .s(n30), .y(\temp[4][29] ) );
  mux21_66 mux21_j_3_6 ( .a(\temp[3][30] ), .b(n17), .s(n30), .y(\temp[4][30] ) );
  mux21_65 mux21_j_3_7 ( .a(\temp[3][31] ), .b(n17), .s(n30), .y(\temp[4][31] ) );
  mux21_64 mux21_k_4_0 ( .a(\temp[4][0] ), .b(\temp[4][16] ), .s(n31), .y(y[0]) );
  mux21_63 mux21_k_4_1 ( .a(\temp[4][1] ), .b(\temp[4][17] ), .s(n31), .y(y[1]) );
  mux21_62 mux21_k_4_2 ( .a(\temp[4][2] ), .b(\temp[4][18] ), .s(n31), .y(y[2]) );
  mux21_61 mux21_k_4_3 ( .a(\temp[4][3] ), .b(\temp[4][19] ), .s(n31), .y(y[3]) );
  mux21_60 mux21_k_4_4 ( .a(\temp[4][4] ), .b(\temp[4][20] ), .s(n31), .y(y[4]) );
  mux21_59 mux21_k_4_5 ( .a(\temp[4][5] ), .b(\temp[4][21] ), .s(n31), .y(y[5]) );
  mux21_58 mux21_k_4_6 ( .a(\temp[4][6] ), .b(\temp[4][22] ), .s(n31), .y(y[6]) );
  mux21_57 mux21_k_4_7 ( .a(\temp[4][7] ), .b(\temp[4][23] ), .s(n31), .y(y[7]) );
  mux21_56 mux21_k_4_8 ( .a(\temp[4][8] ), .b(\temp[4][24] ), .s(n31), .y(y[8]) );
  mux21_55 mux21_k_4_9 ( .a(\temp[4][9] ), .b(\temp[4][25] ), .s(n31), .y(y[9]) );
  mux21_54 mux21_k_4_10 ( .a(\temp[4][10] ), .b(\temp[4][26] ), .s(n31), .y(
        y[10]) );
  mux21_53 mux21_k_4_11 ( .a(\temp[4][11] ), .b(\temp[4][27] ), .s(n31), .y(
        y[11]) );
  mux21_52 mux21_k_4_12 ( .a(\temp[4][12] ), .b(\temp[4][28] ), .s(n32), .y(
        y[12]) );
  mux21_51 mux21_k_4_13 ( .a(\temp[4][13] ), .b(\temp[4][29] ), .s(n32), .y(
        y[13]) );
  mux21_50 mux21_k_4_14 ( .a(\temp[4][14] ), .b(\temp[4][30] ), .s(n32), .y(
        y[14]) );
  mux21_49 mux21_k_4_15 ( .a(\temp[4][15] ), .b(\temp[4][31] ), .s(n32), .y(
        y[15]) );
  mux21_48 mux21_j_4_0 ( .a(\temp[4][16] ), .b(n17), .s(n32), .y(y[16]) );
  mux21_47 mux21_j_4_1 ( .a(\temp[4][17] ), .b(n17), .s(n32), .y(y[17]) );
  mux21_46 mux21_j_4_2 ( .a(\temp[4][18] ), .b(n17), .s(n32), .y(y[18]) );
  mux21_45 mux21_j_4_3 ( .a(\temp[4][19] ), .b(n17), .s(n32), .y(y[19]) );
  mux21_44 mux21_j_4_4 ( .a(\temp[4][20] ), .b(n17), .s(n32), .y(y[20]) );
  mux21_43 mux21_j_4_5 ( .a(\temp[4][21] ), .b(n17), .s(n32), .y(y[21]) );
  mux21_42 mux21_j_4_6 ( .a(\temp[4][22] ), .b(n17), .s(n32), .y(y[22]) );
  mux21_41 mux21_j_4_7 ( .a(\temp[4][23] ), .b(n17), .s(n32), .y(y[23]) );
  mux21_40 mux21_j_4_8 ( .a(\temp[4][24] ), .b(n17), .s(n33), .y(y[24]) );
  mux21_39 mux21_j_4_9 ( .a(\temp[4][25] ), .b(n18), .s(n33), .y(y[25]) );
  mux21_38 mux21_j_4_10 ( .a(\temp[4][26] ), .b(n18), .s(n33), .y(y[26]) );
  mux21_37 mux21_j_4_11 ( .a(\temp[4][27] ), .b(n18), .s(n33), .y(y[27]) );
  mux21_36 mux21_j_4_12 ( .a(\temp[4][28] ), .b(n18), .s(n33), .y(y[28]) );
  mux21_35 mux21_j_4_13 ( .a(\temp[4][29] ), .b(n18), .s(n33), .y(y[29]) );
  mux21_34 mux21_j_4_14 ( .a(\temp[4][30] ), .b(n18), .s(n33), .y(y[30]) );
  mux21_33 mux21_j_4_15 ( .a(\temp[4][31] ), .b(n18), .s(n33), .y(y[31]) );
  BUF_X1 U1 ( .A(n3), .Z(n19) );
  BUF_X1 U2 ( .A(n3), .Z(n20) );
  BUF_X1 U3 ( .A(n6), .Z(n22) );
  BUF_X1 U4 ( .A(n6), .Z(n23) );
  BUF_X1 U5 ( .A(n9), .Z(n26) );
  BUF_X1 U6 ( .A(n3), .Z(n21) );
  BUF_X1 U7 ( .A(n6), .Z(n24) );
  BUF_X1 U8 ( .A(n9), .Z(n25) );
  BUF_X1 U9 ( .A(n12), .Z(n28) );
  BUF_X1 U10 ( .A(n12), .Z(n29) );
  BUF_X1 U11 ( .A(n15), .Z(n31) );
  BUF_X1 U12 ( .A(n15), .Z(n32) );
  BUF_X1 U13 ( .A(n9), .Z(n27) );
  BUF_X1 U14 ( .A(n12), .Z(n30) );
  BUF_X1 U15 ( .A(n15), .Z(n33) );
  BUF_X1 U16 ( .A(shift_type), .Z(n16) );
  BUF_X1 U17 ( .A(shift_type), .Z(n17) );
  BUF_X1 U18 ( .A(shift_type), .Z(n18) );
endmodule


module barrel_shifter_left_n32 ( x, pos, y );
  input [31:0] x;
  input [4:0] pos;
  output [31:0] y;
  wire   \temp[4][31] , \temp[4][30] , \temp[4][29] , \temp[4][28] ,
         \temp[4][27] , \temp[4][26] , \temp[4][25] , \temp[4][24] ,
         \temp[4][23] , \temp[4][22] , \temp[4][21] , \temp[4][20] ,
         \temp[4][19] , \temp[4][18] , \temp[4][17] , \temp[4][16] ,
         \temp[4][15] , \temp[4][14] , \temp[4][13] , \temp[4][12] ,
         \temp[4][11] , \temp[4][10] , \temp[4][9] , \temp[4][8] ,
         \temp[4][7] , \temp[4][6] , \temp[4][5] , \temp[4][4] , \temp[4][3] ,
         \temp[4][2] , \temp[4][1] , \temp[4][0] , \temp[3][31] ,
         \temp[3][30] , \temp[3][29] , \temp[3][28] , \temp[3][27] ,
         \temp[3][26] , \temp[3][25] , \temp[3][24] , \temp[3][23] ,
         \temp[3][22] , \temp[3][21] , \temp[3][20] , \temp[3][19] ,
         \temp[3][18] , \temp[3][17] , \temp[3][16] , \temp[3][15] ,
         \temp[3][14] , \temp[3][13] , \temp[3][12] , \temp[3][11] ,
         \temp[3][10] , \temp[3][9] , \temp[3][8] , \temp[3][7] , \temp[3][6] ,
         \temp[3][5] , \temp[3][4] , \temp[3][3] , \temp[3][2] , \temp[3][1] ,
         \temp[3][0] , \temp[2][31] , \temp[2][30] , \temp[2][29] ,
         \temp[2][28] , \temp[2][27] , \temp[2][26] , \temp[2][25] ,
         \temp[2][24] , \temp[2][23] , \temp[2][22] , \temp[2][21] ,
         \temp[2][20] , \temp[2][19] , \temp[2][18] , \temp[2][17] ,
         \temp[2][16] , \temp[2][15] , \temp[2][14] , \temp[2][13] ,
         \temp[2][12] , \temp[2][11] , \temp[2][10] , \temp[2][9] ,
         \temp[2][8] , \temp[2][7] , \temp[2][6] , \temp[2][5] , \temp[2][4] ,
         \temp[2][3] , \temp[2][2] , \temp[2][1] , \temp[2][0] , \temp[1][31] ,
         \temp[1][30] , \temp[1][29] , \temp[1][28] , \temp[1][27] ,
         \temp[1][26] , \temp[1][25] , \temp[1][24] , \temp[1][23] ,
         \temp[1][22] , \temp[1][21] , \temp[1][20] , \temp[1][19] ,
         \temp[1][18] , \temp[1][17] , \temp[1][16] , \temp[1][15] ,
         \temp[1][14] , \temp[1][13] , \temp[1][12] , \temp[1][11] ,
         \temp[1][10] , \temp[1][9] , \temp[1][8] , \temp[1][7] , \temp[1][6] ,
         \temp[1][5] , \temp[1][4] , \temp[1][3] , \temp[1][2] , \temp[1][1] ,
         \temp[1][0] , n3, n6, n9, n12, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30;
  tri   [31:0] y;
  assign n3 = pos[0];
  assign n6 = pos[1];
  assign n9 = pos[2];
  assign n12 = pos[3];
  assign n15 = pos[4];

  mux21_352 mux21_j_0_0 ( .a(x[0]), .b(1'b0), .s(n16), .y(\temp[1][0] ) );
  mux21_351 mux21_k_0_0 ( .a(x[1]), .b(x[0]), .s(n16), .y(\temp[1][1] ) );
  mux21_350 mux21_k_0_1 ( .a(x[2]), .b(x[1]), .s(n16), .y(\temp[1][2] ) );
  mux21_349 mux21_k_0_2 ( .a(x[3]), .b(x[2]), .s(n16), .y(\temp[1][3] ) );
  mux21_348 mux21_k_0_3 ( .a(x[4]), .b(x[3]), .s(n16), .y(\temp[1][4] ) );
  mux21_347 mux21_k_0_4 ( .a(x[5]), .b(x[4]), .s(n16), .y(\temp[1][5] ) );
  mux21_346 mux21_k_0_5 ( .a(x[6]), .b(x[5]), .s(n16), .y(\temp[1][6] ) );
  mux21_345 mux21_k_0_6 ( .a(x[7]), .b(x[6]), .s(n16), .y(\temp[1][7] ) );
  mux21_344 mux21_k_0_7 ( .a(x[8]), .b(x[7]), .s(n16), .y(\temp[1][8] ) );
  mux21_343 mux21_k_0_8 ( .a(x[9]), .b(x[8]), .s(n16), .y(\temp[1][9] ) );
  mux21_342 mux21_k_0_9 ( .a(x[10]), .b(x[9]), .s(n16), .y(\temp[1][10] ) );
  mux21_341 mux21_k_0_10 ( .a(x[11]), .b(x[10]), .s(n16), .y(\temp[1][11] ) );
  mux21_340 mux21_k_0_11 ( .a(x[12]), .b(x[11]), .s(n17), .y(\temp[1][12] ) );
  mux21_339 mux21_k_0_12 ( .a(x[13]), .b(x[12]), .s(n17), .y(\temp[1][13] ) );
  mux21_338 mux21_k_0_13 ( .a(x[14]), .b(x[13]), .s(n17), .y(\temp[1][14] ) );
  mux21_337 mux21_k_0_14 ( .a(x[15]), .b(x[14]), .s(n17), .y(\temp[1][15] ) );
  mux21_336 mux21_k_0_15 ( .a(x[16]), .b(x[15]), .s(n17), .y(\temp[1][16] ) );
  mux21_335 mux21_k_0_16 ( .a(x[17]), .b(x[16]), .s(n17), .y(\temp[1][17] ) );
  mux21_334 mux21_k_0_17 ( .a(x[18]), .b(x[17]), .s(n17), .y(\temp[1][18] ) );
  mux21_333 mux21_k_0_18 ( .a(x[19]), .b(x[18]), .s(n17), .y(\temp[1][19] ) );
  mux21_332 mux21_k_0_19 ( .a(x[20]), .b(x[19]), .s(n17), .y(\temp[1][20] ) );
  mux21_331 mux21_k_0_20 ( .a(x[21]), .b(x[20]), .s(n17), .y(\temp[1][21] ) );
  mux21_330 mux21_k_0_21 ( .a(x[22]), .b(x[21]), .s(n17), .y(\temp[1][22] ) );
  mux21_329 mux21_k_0_22 ( .a(x[23]), .b(x[22]), .s(n17), .y(\temp[1][23] ) );
  mux21_328 mux21_k_0_23 ( .a(x[24]), .b(x[23]), .s(n18), .y(\temp[1][24] ) );
  mux21_327 mux21_k_0_24 ( .a(x[25]), .b(x[24]), .s(n18), .y(\temp[1][25] ) );
  mux21_326 mux21_k_0_25 ( .a(x[26]), .b(x[25]), .s(n18), .y(\temp[1][26] ) );
  mux21_325 mux21_k_0_26 ( .a(x[27]), .b(x[26]), .s(n18), .y(\temp[1][27] ) );
  mux21_324 mux21_k_0_27 ( .a(x[28]), .b(x[27]), .s(n18), .y(\temp[1][28] ) );
  mux21_323 mux21_k_0_28 ( .a(x[29]), .b(x[28]), .s(n18), .y(\temp[1][29] ) );
  mux21_322 mux21_k_0_29 ( .a(x[30]), .b(x[29]), .s(n18), .y(\temp[1][30] ) );
  mux21_321 mux21_k_0_30 ( .a(x[31]), .b(x[30]), .s(n18), .y(\temp[1][31] ) );
  mux21_320 mux21_j_1_0 ( .a(\temp[1][0] ), .b(1'b0), .s(n19), .y(\temp[2][0] ) );
  mux21_319 mux21_j_1_1 ( .a(\temp[1][1] ), .b(1'b0), .s(n19), .y(\temp[2][1] ) );
  mux21_318 mux21_k_1_0 ( .a(\temp[1][2] ), .b(\temp[1][0] ), .s(n19), .y(
        \temp[2][2] ) );
  mux21_317 mux21_k_1_1 ( .a(\temp[1][3] ), .b(\temp[1][1] ), .s(n19), .y(
        \temp[2][3] ) );
  mux21_316 mux21_k_1_2 ( .a(\temp[1][4] ), .b(\temp[1][2] ), .s(n19), .y(
        \temp[2][4] ) );
  mux21_315 mux21_k_1_3 ( .a(\temp[1][5] ), .b(\temp[1][3] ), .s(n19), .y(
        \temp[2][5] ) );
  mux21_314 mux21_k_1_4 ( .a(\temp[1][6] ), .b(\temp[1][4] ), .s(n19), .y(
        \temp[2][6] ) );
  mux21_313 mux21_k_1_5 ( .a(\temp[1][7] ), .b(\temp[1][5] ), .s(n19), .y(
        \temp[2][7] ) );
  mux21_312 mux21_k_1_6 ( .a(\temp[1][8] ), .b(\temp[1][6] ), .s(n19), .y(
        \temp[2][8] ) );
  mux21_311 mux21_k_1_7 ( .a(\temp[1][9] ), .b(\temp[1][7] ), .s(n19), .y(
        \temp[2][9] ) );
  mux21_310 mux21_k_1_8 ( .a(\temp[1][10] ), .b(\temp[1][8] ), .s(n19), .y(
        \temp[2][10] ) );
  mux21_309 mux21_k_1_9 ( .a(\temp[1][11] ), .b(\temp[1][9] ), .s(n19), .y(
        \temp[2][11] ) );
  mux21_308 mux21_k_1_10 ( .a(\temp[1][12] ), .b(\temp[1][10] ), .s(n20), .y(
        \temp[2][12] ) );
  mux21_307 mux21_k_1_11 ( .a(\temp[1][13] ), .b(\temp[1][11] ), .s(n20), .y(
        \temp[2][13] ) );
  mux21_306 mux21_k_1_12 ( .a(\temp[1][14] ), .b(\temp[1][12] ), .s(n20), .y(
        \temp[2][14] ) );
  mux21_305 mux21_k_1_13 ( .a(\temp[1][15] ), .b(\temp[1][13] ), .s(n20), .y(
        \temp[2][15] ) );
  mux21_304 mux21_k_1_14 ( .a(\temp[1][16] ), .b(\temp[1][14] ), .s(n20), .y(
        \temp[2][16] ) );
  mux21_303 mux21_k_1_15 ( .a(\temp[1][17] ), .b(\temp[1][15] ), .s(n20), .y(
        \temp[2][17] ) );
  mux21_302 mux21_k_1_16 ( .a(\temp[1][18] ), .b(\temp[1][16] ), .s(n20), .y(
        \temp[2][18] ) );
  mux21_301 mux21_k_1_17 ( .a(\temp[1][19] ), .b(\temp[1][17] ), .s(n20), .y(
        \temp[2][19] ) );
  mux21_300 mux21_k_1_18 ( .a(\temp[1][20] ), .b(\temp[1][18] ), .s(n20), .y(
        \temp[2][20] ) );
  mux21_299 mux21_k_1_19 ( .a(\temp[1][21] ), .b(\temp[1][19] ), .s(n20), .y(
        \temp[2][21] ) );
  mux21_298 mux21_k_1_20 ( .a(\temp[1][22] ), .b(\temp[1][20] ), .s(n20), .y(
        \temp[2][22] ) );
  mux21_297 mux21_k_1_21 ( .a(\temp[1][23] ), .b(\temp[1][21] ), .s(n20), .y(
        \temp[2][23] ) );
  mux21_296 mux21_k_1_22 ( .a(\temp[1][24] ), .b(\temp[1][22] ), .s(n21), .y(
        \temp[2][24] ) );
  mux21_295 mux21_k_1_23 ( .a(\temp[1][25] ), .b(\temp[1][23] ), .s(n21), .y(
        \temp[2][25] ) );
  mux21_294 mux21_k_1_24 ( .a(\temp[1][26] ), .b(\temp[1][24] ), .s(n21), .y(
        \temp[2][26] ) );
  mux21_293 mux21_k_1_25 ( .a(\temp[1][27] ), .b(\temp[1][25] ), .s(n21), .y(
        \temp[2][27] ) );
  mux21_292 mux21_k_1_26 ( .a(\temp[1][28] ), .b(\temp[1][26] ), .s(n21), .y(
        \temp[2][28] ) );
  mux21_291 mux21_k_1_27 ( .a(\temp[1][29] ), .b(\temp[1][27] ), .s(n21), .y(
        \temp[2][29] ) );
  mux21_290 mux21_k_1_28 ( .a(\temp[1][30] ), .b(\temp[1][28] ), .s(n21), .y(
        \temp[2][30] ) );
  mux21_289 mux21_k_1_29 ( .a(\temp[1][31] ), .b(\temp[1][29] ), .s(n21), .y(
        \temp[2][31] ) );
  mux21_288 mux21_j_2_0 ( .a(\temp[2][0] ), .b(1'b0), .s(n22), .y(\temp[3][0] ) );
  mux21_287 mux21_j_2_1 ( .a(\temp[2][1] ), .b(1'b0), .s(n22), .y(\temp[3][1] ) );
  mux21_286 mux21_j_2_2 ( .a(\temp[2][2] ), .b(1'b0), .s(n22), .y(\temp[3][2] ) );
  mux21_285 mux21_j_2_3 ( .a(\temp[2][3] ), .b(1'b0), .s(n22), .y(\temp[3][3] ) );
  mux21_284 mux21_k_2_0 ( .a(\temp[2][4] ), .b(\temp[2][0] ), .s(n22), .y(
        \temp[3][4] ) );
  mux21_283 mux21_k_2_1 ( .a(\temp[2][5] ), .b(\temp[2][1] ), .s(n22), .y(
        \temp[3][5] ) );
  mux21_282 mux21_k_2_2 ( .a(\temp[2][6] ), .b(\temp[2][2] ), .s(n22), .y(
        \temp[3][6] ) );
  mux21_281 mux21_k_2_3 ( .a(\temp[2][7] ), .b(\temp[2][3] ), .s(n22), .y(
        \temp[3][7] ) );
  mux21_280 mux21_k_2_4 ( .a(\temp[2][8] ), .b(\temp[2][4] ), .s(n22), .y(
        \temp[3][8] ) );
  mux21_279 mux21_k_2_5 ( .a(\temp[2][9] ), .b(\temp[2][5] ), .s(n22), .y(
        \temp[3][9] ) );
  mux21_278 mux21_k_2_6 ( .a(\temp[2][10] ), .b(\temp[2][6] ), .s(n22), .y(
        \temp[3][10] ) );
  mux21_277 mux21_k_2_7 ( .a(\temp[2][11] ), .b(\temp[2][7] ), .s(n22), .y(
        \temp[3][11] ) );
  mux21_276 mux21_k_2_8 ( .a(\temp[2][12] ), .b(\temp[2][8] ), .s(n23), .y(
        \temp[3][12] ) );
  mux21_275 mux21_k_2_9 ( .a(\temp[2][13] ), .b(\temp[2][9] ), .s(n23), .y(
        \temp[3][13] ) );
  mux21_274 mux21_k_2_10 ( .a(\temp[2][14] ), .b(\temp[2][10] ), .s(n23), .y(
        \temp[3][14] ) );
  mux21_273 mux21_k_2_11 ( .a(\temp[2][15] ), .b(\temp[2][11] ), .s(n23), .y(
        \temp[3][15] ) );
  mux21_272 mux21_k_2_12 ( .a(\temp[2][16] ), .b(\temp[2][12] ), .s(n23), .y(
        \temp[3][16] ) );
  mux21_271 mux21_k_2_13 ( .a(\temp[2][17] ), .b(\temp[2][13] ), .s(n23), .y(
        \temp[3][17] ) );
  mux21_270 mux21_k_2_14 ( .a(\temp[2][18] ), .b(\temp[2][14] ), .s(n23), .y(
        \temp[3][18] ) );
  mux21_269 mux21_k_2_15 ( .a(\temp[2][19] ), .b(\temp[2][15] ), .s(n23), .y(
        \temp[3][19] ) );
  mux21_268 mux21_k_2_16 ( .a(\temp[2][20] ), .b(\temp[2][16] ), .s(n23), .y(
        \temp[3][20] ) );
  mux21_267 mux21_k_2_17 ( .a(\temp[2][21] ), .b(\temp[2][17] ), .s(n23), .y(
        \temp[3][21] ) );
  mux21_266 mux21_k_2_18 ( .a(\temp[2][22] ), .b(\temp[2][18] ), .s(n23), .y(
        \temp[3][22] ) );
  mux21_265 mux21_k_2_19 ( .a(\temp[2][23] ), .b(\temp[2][19] ), .s(n23), .y(
        \temp[3][23] ) );
  mux21_264 mux21_k_2_20 ( .a(\temp[2][24] ), .b(\temp[2][20] ), .s(n24), .y(
        \temp[3][24] ) );
  mux21_263 mux21_k_2_21 ( .a(\temp[2][25] ), .b(\temp[2][21] ), .s(n24), .y(
        \temp[3][25] ) );
  mux21_262 mux21_k_2_22 ( .a(\temp[2][26] ), .b(\temp[2][22] ), .s(n24), .y(
        \temp[3][26] ) );
  mux21_261 mux21_k_2_23 ( .a(\temp[2][27] ), .b(\temp[2][23] ), .s(n24), .y(
        \temp[3][27] ) );
  mux21_260 mux21_k_2_24 ( .a(\temp[2][28] ), .b(\temp[2][24] ), .s(n24), .y(
        \temp[3][28] ) );
  mux21_259 mux21_k_2_25 ( .a(\temp[2][29] ), .b(\temp[2][25] ), .s(n24), .y(
        \temp[3][29] ) );
  mux21_258 mux21_k_2_26 ( .a(\temp[2][30] ), .b(\temp[2][26] ), .s(n24), .y(
        \temp[3][30] ) );
  mux21_257 mux21_k_2_27 ( .a(\temp[2][31] ), .b(\temp[2][27] ), .s(n24), .y(
        \temp[3][31] ) );
  mux21_256 mux21_j_3_0 ( .a(\temp[3][0] ), .b(1'b0), .s(n25), .y(\temp[4][0] ) );
  mux21_255 mux21_j_3_1 ( .a(\temp[3][1] ), .b(1'b0), .s(n25), .y(\temp[4][1] ) );
  mux21_254 mux21_j_3_2 ( .a(\temp[3][2] ), .b(1'b0), .s(n25), .y(\temp[4][2] ) );
  mux21_253 mux21_j_3_3 ( .a(\temp[3][3] ), .b(1'b0), .s(n25), .y(\temp[4][3] ) );
  mux21_252 mux21_j_3_4 ( .a(\temp[3][4] ), .b(1'b0), .s(n25), .y(\temp[4][4] ) );
  mux21_251 mux21_j_3_5 ( .a(\temp[3][5] ), .b(1'b0), .s(n25), .y(\temp[4][5] ) );
  mux21_250 mux21_j_3_6 ( .a(\temp[3][6] ), .b(1'b0), .s(n25), .y(\temp[4][6] ) );
  mux21_249 mux21_j_3_7 ( .a(\temp[3][7] ), .b(1'b0), .s(n25), .y(\temp[4][7] ) );
  mux21_248 mux21_k_3_0 ( .a(\temp[3][8] ), .b(\temp[3][0] ), .s(n25), .y(
        \temp[4][8] ) );
  mux21_247 mux21_k_3_1 ( .a(\temp[3][9] ), .b(\temp[3][1] ), .s(n25), .y(
        \temp[4][9] ) );
  mux21_246 mux21_k_3_2 ( .a(\temp[3][10] ), .b(\temp[3][2] ), .s(n25), .y(
        \temp[4][10] ) );
  mux21_245 mux21_k_3_3 ( .a(\temp[3][11] ), .b(\temp[3][3] ), .s(n25), .y(
        \temp[4][11] ) );
  mux21_244 mux21_k_3_4 ( .a(\temp[3][12] ), .b(\temp[3][4] ), .s(n26), .y(
        \temp[4][12] ) );
  mux21_243 mux21_k_3_5 ( .a(\temp[3][13] ), .b(\temp[3][5] ), .s(n26), .y(
        \temp[4][13] ) );
  mux21_242 mux21_k_3_6 ( .a(\temp[3][14] ), .b(\temp[3][6] ), .s(n26), .y(
        \temp[4][14] ) );
  mux21_241 mux21_k_3_7 ( .a(\temp[3][15] ), .b(\temp[3][7] ), .s(n26), .y(
        \temp[4][15] ) );
  mux21_240 mux21_k_3_8 ( .a(\temp[3][16] ), .b(\temp[3][8] ), .s(n26), .y(
        \temp[4][16] ) );
  mux21_239 mux21_k_3_9 ( .a(\temp[3][17] ), .b(\temp[3][9] ), .s(n26), .y(
        \temp[4][17] ) );
  mux21_238 mux21_k_3_10 ( .a(\temp[3][18] ), .b(\temp[3][10] ), .s(n26), .y(
        \temp[4][18] ) );
  mux21_237 mux21_k_3_11 ( .a(\temp[3][19] ), .b(\temp[3][11] ), .s(n26), .y(
        \temp[4][19] ) );
  mux21_236 mux21_k_3_12 ( .a(\temp[3][20] ), .b(\temp[3][12] ), .s(n26), .y(
        \temp[4][20] ) );
  mux21_235 mux21_k_3_13 ( .a(\temp[3][21] ), .b(\temp[3][13] ), .s(n26), .y(
        \temp[4][21] ) );
  mux21_234 mux21_k_3_14 ( .a(\temp[3][22] ), .b(\temp[3][14] ), .s(n26), .y(
        \temp[4][22] ) );
  mux21_233 mux21_k_3_15 ( .a(\temp[3][23] ), .b(\temp[3][15] ), .s(n26), .y(
        \temp[4][23] ) );
  mux21_232 mux21_k_3_16 ( .a(\temp[3][24] ), .b(\temp[3][16] ), .s(n27), .y(
        \temp[4][24] ) );
  mux21_231 mux21_k_3_17 ( .a(\temp[3][25] ), .b(\temp[3][17] ), .s(n27), .y(
        \temp[4][25] ) );
  mux21_230 mux21_k_3_18 ( .a(\temp[3][26] ), .b(\temp[3][18] ), .s(n27), .y(
        \temp[4][26] ) );
  mux21_229 mux21_k_3_19 ( .a(\temp[3][27] ), .b(\temp[3][19] ), .s(n27), .y(
        \temp[4][27] ) );
  mux21_228 mux21_k_3_20 ( .a(\temp[3][28] ), .b(\temp[3][20] ), .s(n27), .y(
        \temp[4][28] ) );
  mux21_227 mux21_k_3_21 ( .a(\temp[3][29] ), .b(\temp[3][21] ), .s(n27), .y(
        \temp[4][29] ) );
  mux21_226 mux21_k_3_22 ( .a(\temp[3][30] ), .b(\temp[3][22] ), .s(n27), .y(
        \temp[4][30] ) );
  mux21_225 mux21_k_3_23 ( .a(\temp[3][31] ), .b(\temp[3][23] ), .s(n27), .y(
        \temp[4][31] ) );
  mux21_224 mux21_j_4_0 ( .a(\temp[4][0] ), .b(1'b0), .s(n28), .y(y[0]) );
  mux21_223 mux21_j_4_1 ( .a(\temp[4][1] ), .b(1'b0), .s(n28), .y(y[1]) );
  mux21_222 mux21_j_4_2 ( .a(\temp[4][2] ), .b(1'b0), .s(n28), .y(y[2]) );
  mux21_221 mux21_j_4_3 ( .a(\temp[4][3] ), .b(1'b0), .s(n28), .y(y[3]) );
  mux21_220 mux21_j_4_4 ( .a(\temp[4][4] ), .b(1'b0), .s(n28), .y(y[4]) );
  mux21_219 mux21_j_4_5 ( .a(\temp[4][5] ), .b(1'b0), .s(n28), .y(y[5]) );
  mux21_218 mux21_j_4_6 ( .a(\temp[4][6] ), .b(1'b0), .s(n28), .y(y[6]) );
  mux21_217 mux21_j_4_7 ( .a(\temp[4][7] ), .b(1'b0), .s(n28), .y(y[7]) );
  mux21_216 mux21_j_4_8 ( .a(\temp[4][8] ), .b(1'b0), .s(n28), .y(y[8]) );
  mux21_215 mux21_j_4_9 ( .a(\temp[4][9] ), .b(1'b0), .s(n28), .y(y[9]) );
  mux21_214 mux21_j_4_10 ( .a(\temp[4][10] ), .b(1'b0), .s(n28), .y(y[10]) );
  mux21_213 mux21_j_4_11 ( .a(\temp[4][11] ), .b(1'b0), .s(n28), .y(y[11]) );
  mux21_212 mux21_j_4_12 ( .a(\temp[4][12] ), .b(1'b0), .s(n29), .y(y[12]) );
  mux21_211 mux21_j_4_13 ( .a(\temp[4][13] ), .b(1'b0), .s(n29), .y(y[13]) );
  mux21_210 mux21_j_4_14 ( .a(\temp[4][14] ), .b(1'b0), .s(n29), .y(y[14]) );
  mux21_209 mux21_j_4_15 ( .a(\temp[4][15] ), .b(1'b0), .s(n29), .y(y[15]) );
  mux21_208 mux21_k_4_0 ( .a(\temp[4][16] ), .b(\temp[4][0] ), .s(n29), .y(
        y[16]) );
  mux21_207 mux21_k_4_1 ( .a(\temp[4][17] ), .b(\temp[4][1] ), .s(n29), .y(
        y[17]) );
  mux21_206 mux21_k_4_2 ( .a(\temp[4][18] ), .b(\temp[4][2] ), .s(n29), .y(
        y[18]) );
  mux21_205 mux21_k_4_3 ( .a(\temp[4][19] ), .b(\temp[4][3] ), .s(n29), .y(
        y[19]) );
  mux21_204 mux21_k_4_4 ( .a(\temp[4][20] ), .b(\temp[4][4] ), .s(n29), .y(
        y[20]) );
  mux21_203 mux21_k_4_5 ( .a(\temp[4][21] ), .b(\temp[4][5] ), .s(n29), .y(
        y[21]) );
  mux21_202 mux21_k_4_6 ( .a(\temp[4][22] ), .b(\temp[4][6] ), .s(n29), .y(
        y[22]) );
  mux21_201 mux21_k_4_7 ( .a(\temp[4][23] ), .b(\temp[4][7] ), .s(n29), .y(
        y[23]) );
  mux21_200 mux21_k_4_8 ( .a(\temp[4][24] ), .b(\temp[4][8] ), .s(n30), .y(
        y[24]) );
  mux21_199 mux21_k_4_9 ( .a(\temp[4][25] ), .b(\temp[4][9] ), .s(n30), .y(
        y[25]) );
  mux21_198 mux21_k_4_10 ( .a(\temp[4][26] ), .b(\temp[4][10] ), .s(n30), .y(
        y[26]) );
  mux21_197 mux21_k_4_11 ( .a(\temp[4][27] ), .b(\temp[4][11] ), .s(n30), .y(
        y[27]) );
  mux21_196 mux21_k_4_12 ( .a(\temp[4][28] ), .b(\temp[4][12] ), .s(n30), .y(
        y[28]) );
  mux21_195 mux21_k_4_13 ( .a(\temp[4][29] ), .b(\temp[4][13] ), .s(n30), .y(
        y[29]) );
  mux21_194 mux21_k_4_14 ( .a(\temp[4][30] ), .b(\temp[4][14] ), .s(n30), .y(
        y[30]) );
  mux21_193 mux21_k_4_15 ( .a(\temp[4][31] ), .b(\temp[4][15] ), .s(n30), .y(
        y[31]) );
  BUF_X1 U2 ( .A(n3), .Z(n17) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  BUF_X1 U4 ( .A(n6), .Z(n20) );
  BUF_X1 U5 ( .A(n6), .Z(n19) );
  BUF_X1 U6 ( .A(n9), .Z(n23) );
  BUF_X1 U7 ( .A(n9), .Z(n22) );
  BUF_X1 U8 ( .A(n3), .Z(n18) );
  BUF_X1 U9 ( .A(n6), .Z(n21) );
  BUF_X1 U10 ( .A(n12), .Z(n25) );
  BUF_X1 U11 ( .A(n12), .Z(n26) );
  BUF_X1 U12 ( .A(n15), .Z(n28) );
  BUF_X1 U13 ( .A(n15), .Z(n29) );
  BUF_X1 U14 ( .A(n9), .Z(n24) );
  BUF_X1 U15 ( .A(n12), .Z(n27) );
  BUF_X1 U16 ( .A(n15), .Z(n30) );
endmodule


module subtractor_n32 ( a, b, cin, y, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input cin;
  output cout;

  wire   [31:0] b_not;

  not_n_n32_0 inv ( .a(b), .y(b_not) );
  rca_n_n32_2 sub ( .a(a), .b(b_not), .c_in(1'b1), .sum(y), .c_out(cout) );
endmodule


module p4_n32 ( a, b, cin, s, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] s;
  input cin;
  output cout;

  wire   [31:0] c_p4;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23;

  sparse_tree_carry_gen_n32 sparse_tree_carry_gen_p4 ( .a(a), .b(b), .c({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, c_p4[7:0]}) );
  sum_generator_n32 sum_generator_p4 ( .a(a), .b(b), .c({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, c_p4[7:0]}), 
        .cin(cin), .s(s), .cout(cout) );
endmodule


module mux21_0 ( a, b, s, y );
  input a, b, s;
  output y;
  wire   sa, y1, y2;

  not_1_0 inv ( .a(s), .y(sa) );
  and_2_1311 and1 ( .a(a), .b(sa), .y(y1) );
  and_2_1310 and2 ( .a(b), .b(s), .y(y2) );
  or_2_644 or1 ( .a(y1), .b(y2), .y(y) );
endmodule


module and_n1_n32 ( a, y );
  input [31:0] a;
  output y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR4_X1 U1 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NAND4_X1 U2 ( .A1(a[12]), .A2(a[11]), .A3(a[10]), .A4(a[0]), .ZN(n3) );
  NAND4_X1 U3 ( .A1(a[16]), .A2(a[15]), .A3(a[14]), .A4(a[13]), .ZN(n4) );
  NAND4_X1 U4 ( .A1(a[1]), .A2(a[19]), .A3(a[18]), .A4(a[17]), .ZN(n5) );
  AND2_X1 U5 ( .A1(n1), .A2(n2), .ZN(y) );
  NOR4_X1 U6 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NAND4_X1 U7 ( .A1(a[23]), .A2(a[22]), .A3(a[21]), .A4(a[20]), .ZN(n6) );
  NAND4_X1 U8 ( .A1(a[9]), .A2(a[8]), .A3(a[7]), .A4(a[6]), .ZN(n10) );
  NAND4_X1 U9 ( .A1(a[5]), .A2(a[4]), .A3(a[3]), .A4(a[31]), .ZN(n9) );
  NAND4_X1 U10 ( .A1(a[30]), .A2(a[2]), .A3(a[29]), .A4(a[28]), .ZN(n8) );
  NAND4_X1 U11 ( .A1(a[27]), .A2(a[26]), .A3(a[25]), .A4(a[24]), .ZN(n7) );
endmodule


module xnor_2_0 ( a, b, y );
  input a, b;
  output y;


  XNOR2_X1 U1 ( .A(b), .B(a), .ZN(y) );
endmodule


module fa_2_0 ( a, b, c_in, sum, c_out );
  input a, b, c_in;
  output sum, c_out;
  wire   s1, s3, s2;

  xor_2_352 xor1 ( .a(a), .b(b), .y(s1) );
  xor_2_351 xor2 ( .a(s1), .b(c_in), .y(sum) );
  and_2_1375 and1 ( .a(a), .b(b), .y(s3) );
  and_2_1374 and2 ( .a(s1), .b(c_in), .y(s2) );
  or_2_0 or1 ( .a(s2), .b(s3), .y(c_out) );
endmodule


module ffd_async_289 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module ffd_async_291 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;
  wire   n1;

  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q), .QN(n1) );
endmodule


module ffd_async_0 ( clk, reset, en, d, q );
  input clk, reset, en, d;
  output q;


  DFFR_X1 q_reg ( .D(d), .CK(clk), .RN(reset), .Q(q) );
endmodule


module alu_nbit32 ( a, b, unit_sel, y );
  input [31:0] a;
  input [31:0] b;
  input [3:0] unit_sel;
  output [31:0] y;
  wire   type_sr, \cmp_out[0] , \eq_out[0] ;
  wire   [31:0] out_add;
  wire   [31:0] out_sub;
  wire   [31:0] out_log;
  tri   [31:0] out_sl;

  p4_n32 add ( .a(a), .b(b), .cin(1'b0), .s(out_add) );
  subtractor_n32 sub ( .a(a), .b(b), .cin(1'b0), .y(out_sub) );
  barrel_shifter_left_n32 sl ( .x(a), .pos(b[4:0]), .y(out_sl) );
  barrel_shifter_right_n32 sr ( .x(a), .pos(b[4:0]), .shift_type(type_sr), .y(
        out_sl) );
  comparator_n32 comp ( .a(a), .b(b), .cout(\cmp_out[0] ), .z(\eq_out[0] ) );
  xor_2_353 sh ( .a(unit_sel[2]), .b(unit_sel[0]), .y(type_sr) );
  logic_n_n32 logi ( .r1(a), .r2(b), .s0(unit_sel[0]), .s1(unit_sel[1]), .s2(
        unit_sel[2]), .s3(unit_sel[3]), .y(out_log) );
  encoder_n32 enc ( .out_add(out_add), .out_sub(out_sub), .out_sl(out_sl), 
        .out_sr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .out_log(out_log), .out_cmp({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \cmp_out[0] }), .out_eq({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \eq_out[0] }), .sel(unit_sel), .o(y) );
endmodule


module mux21_generic_n32_0 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n1, n2, n3;

  mux21_0 mux21_i_0 ( .a(a[0]), .b(b[0]), .s(n3), .y(y[0]) );
  mux21_479 mux21_i_1 ( .a(a[1]), .b(b[1]), .s(n1), .y(y[1]) );
  mux21_478 mux21_i_2 ( .a(a[2]), .b(b[2]), .s(n1), .y(y[2]) );
  mux21_477 mux21_i_3 ( .a(a[3]), .b(b[3]), .s(n1), .y(y[3]) );
  mux21_476 mux21_i_4 ( .a(a[4]), .b(b[4]), .s(n1), .y(y[4]) );
  mux21_475 mux21_i_5 ( .a(a[5]), .b(b[5]), .s(n1), .y(y[5]) );
  mux21_474 mux21_i_6 ( .a(a[6]), .b(b[6]), .s(n1), .y(y[6]) );
  mux21_473 mux21_i_7 ( .a(a[7]), .b(b[7]), .s(n1), .y(y[7]) );
  mux21_472 mux21_i_8 ( .a(a[8]), .b(b[8]), .s(n1), .y(y[8]) );
  mux21_471 mux21_i_9 ( .a(a[9]), .b(b[9]), .s(n1), .y(y[9]) );
  mux21_470 mux21_i_10 ( .a(a[10]), .b(b[10]), .s(n1), .y(y[10]) );
  mux21_469 mux21_i_11 ( .a(a[11]), .b(b[11]), .s(n1), .y(y[11]) );
  mux21_468 mux21_i_12 ( .a(a[12]), .b(b[12]), .s(n1), .y(y[12]) );
  mux21_467 mux21_i_13 ( .a(a[13]), .b(b[13]), .s(n2), .y(y[13]) );
  mux21_466 mux21_i_14 ( .a(a[14]), .b(b[14]), .s(n2), .y(y[14]) );
  mux21_465 mux21_i_15 ( .a(a[15]), .b(b[15]), .s(n2), .y(y[15]) );
  mux21_464 mux21_i_16 ( .a(a[16]), .b(b[16]), .s(n2), .y(y[16]) );
  mux21_463 mux21_i_17 ( .a(a[17]), .b(b[17]), .s(n2), .y(y[17]) );
  mux21_462 mux21_i_18 ( .a(a[18]), .b(b[18]), .s(n2), .y(y[18]) );
  mux21_461 mux21_i_19 ( .a(a[19]), .b(b[19]), .s(n2), .y(y[19]) );
  mux21_460 mux21_i_20 ( .a(a[20]), .b(b[20]), .s(n2), .y(y[20]) );
  mux21_459 mux21_i_21 ( .a(a[21]), .b(b[21]), .s(n2), .y(y[21]) );
  mux21_458 mux21_i_22 ( .a(a[22]), .b(b[22]), .s(n2), .y(y[22]) );
  mux21_457 mux21_i_23 ( .a(a[23]), .b(b[23]), .s(n2), .y(y[23]) );
  mux21_456 mux21_i_24 ( .a(a[24]), .b(b[24]), .s(n2), .y(y[24]) );
  mux21_455 mux21_i_25 ( .a(a[25]), .b(b[25]), .s(n3), .y(y[25]) );
  mux21_454 mux21_i_26 ( .a(a[26]), .b(b[26]), .s(n3), .y(y[26]) );
  mux21_453 mux21_i_27 ( .a(a[27]), .b(b[27]), .s(n3), .y(y[27]) );
  mux21_452 mux21_i_28 ( .a(a[28]), .b(b[28]), .s(n3), .y(y[28]) );
  mux21_451 mux21_i_29 ( .a(a[29]), .b(b[29]), .s(n3), .y(y[29]) );
  mux21_450 mux21_i_30 ( .a(a[30]), .b(b[30]), .s(n3), .y(y[30]) );
  mux21_449 mux21_i_31 ( .a(a[31]), .b(b[31]), .s(n3), .y(y[31]) );
  BUF_X1 U1 ( .A(sel), .Z(n1) );
  BUF_X1 U2 ( .A(sel), .Z(n3) );
  BUF_X1 U3 ( .A(sel), .Z(n2) );
endmodule


module and_2_0 ( a, b, y );
  input a, b;
  output y;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(y) );
endmodule


module xor_2_0 ( a, b, y );
  input a, b;
  output y;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(y) );
endmodule


module zero_comp_n32 ( x, y );
  input [31:0] x;
  output y;

  wire   [31:0] res;

  xnor_2_0 xnor_i_0 ( .a(x[0]), .b(1'b0), .y(res[0]) );
  xnor_2_31 xnor_i_1 ( .a(x[1]), .b(1'b0), .y(res[1]) );
  xnor_2_30 xnor_i_2 ( .a(x[2]), .b(1'b0), .y(res[2]) );
  xnor_2_29 xnor_i_3 ( .a(x[3]), .b(1'b0), .y(res[3]) );
  xnor_2_28 xnor_i_4 ( .a(x[4]), .b(1'b0), .y(res[4]) );
  xnor_2_27 xnor_i_5 ( .a(x[5]), .b(1'b0), .y(res[5]) );
  xnor_2_26 xnor_i_6 ( .a(x[6]), .b(1'b0), .y(res[6]) );
  xnor_2_25 xnor_i_7 ( .a(x[7]), .b(1'b0), .y(res[7]) );
  xnor_2_24 xnor_i_8 ( .a(x[8]), .b(1'b0), .y(res[8]) );
  xnor_2_23 xnor_i_9 ( .a(x[9]), .b(1'b0), .y(res[9]) );
  xnor_2_22 xnor_i_10 ( .a(x[10]), .b(1'b0), .y(res[10]) );
  xnor_2_21 xnor_i_11 ( .a(x[11]), .b(1'b0), .y(res[11]) );
  xnor_2_20 xnor_i_12 ( .a(x[12]), .b(1'b0), .y(res[12]) );
  xnor_2_19 xnor_i_13 ( .a(x[13]), .b(1'b0), .y(res[13]) );
  xnor_2_18 xnor_i_14 ( .a(x[14]), .b(1'b0), .y(res[14]) );
  xnor_2_17 xnor_i_15 ( .a(x[15]), .b(1'b0), .y(res[15]) );
  xnor_2_16 xnor_i_16 ( .a(x[16]), .b(1'b0), .y(res[16]) );
  xnor_2_15 xnor_i_17 ( .a(x[17]), .b(1'b0), .y(res[17]) );
  xnor_2_14 xnor_i_18 ( .a(x[18]), .b(1'b0), .y(res[18]) );
  xnor_2_13 xnor_i_19 ( .a(x[19]), .b(1'b0), .y(res[19]) );
  xnor_2_12 xnor_i_20 ( .a(x[20]), .b(1'b0), .y(res[20]) );
  xnor_2_11 xnor_i_21 ( .a(x[21]), .b(1'b0), .y(res[21]) );
  xnor_2_10 xnor_i_22 ( .a(x[22]), .b(1'b0), .y(res[22]) );
  xnor_2_9 xnor_i_23 ( .a(x[23]), .b(1'b0), .y(res[23]) );
  xnor_2_8 xnor_i_24 ( .a(x[24]), .b(1'b0), .y(res[24]) );
  xnor_2_7 xnor_i_25 ( .a(x[25]), .b(1'b0), .y(res[25]) );
  xnor_2_6 xnor_i_26 ( .a(x[26]), .b(1'b0), .y(res[26]) );
  xnor_2_5 xnor_i_27 ( .a(x[27]), .b(1'b0), .y(res[27]) );
  xnor_2_4 xnor_i_28 ( .a(x[28]), .b(1'b0), .y(res[28]) );
  xnor_2_3 xnor_i_29 ( .a(x[29]), .b(1'b0), .y(res[29]) );
  xnor_2_2 xnor_i_30 ( .a(x[30]), .b(1'b0), .y(res[30]) );
  xnor_2_1 xnor_i_31 ( .a(x[31]), .b(1'b0), .y(res[31]) );
  and_n1_n32 big_and ( .a(res), .y(y) );
endmodule


module reg_n_n5_0 ( clock, reset, enable, x, y );
  input [4:0] x;
  output [4:0] y;
  input clock, reset, enable;


  ffd_async_143 ff_0 ( .clk(clock), .reset(reset), .en(enable), .d(x[0]), .q(
        y[0]) );
  ffd_async_142 ff_1 ( .clk(clock), .reset(reset), .en(enable), .d(x[1]), .q(
        y[1]) );
  ffd_async_141 ff_2 ( .clk(clock), .reset(reset), .en(enable), .d(x[2]), .q(
        y[2]) );
  ffd_async_140 ff_3 ( .clk(clock), .reset(reset), .en(enable), .d(x[3]), .q(
        y[3]) );
  ffd_async_139 ff_4 ( .clk(clock), .reset(reset), .en(enable), .d(x[4]), .q(
        y[4]) );
endmodule


module sign_extension_s16_f32 ( x, y );
  input [15:0] x;
  output [31:0] y;

  assign y[31] = x[15];
  assign y[30] = x[15];
  assign y[29] = x[15];
  assign y[28] = x[15];
  assign y[27] = x[15];
  assign y[26] = x[15];
  assign y[25] = x[15];
  assign y[24] = x[15];
  assign y[23] = x[15];
  assign y[22] = x[15];
  assign y[21] = x[15];
  assign y[20] = x[15];
  assign y[19] = x[15];
  assign y[18] = x[15];
  assign y[17] = x[15];
  assign y[16] = x[15];
  assign y[15] = x[15];
  assign y[14] = x[14];
  assign y[13] = x[13];
  assign y[12] = x[12];
  assign y[11] = x[11];
  assign y[10] = x[10];
  assign y[9] = x[9];
  assign y[8] = x[8];
  assign y[7] = x[7];
  assign y[6] = x[6];
  assign y[5] = x[5];
  assign y[4] = x[4];
  assign y[3] = x[3];
  assign y[2] = x[2];
  assign y[1] = x[1];
  assign y[0] = x[0];

endmodule


module register_file_n32 ( clk, reset, enable, rd1, rd2, wr, add_wr, add_rd1, 
        add_rd2, datain, out1, out2 );
  input [4:0] add_wr;
  input [4:0] add_rd1;
  input [4:0] add_rd2;
  input [31:0] datain;
  output [31:0] out1;
  output [31:0] out2;
  input clk, reset, enable, rd1, rd2, wr;
  wire   \registers[0][31] , \registers[0][30] , \registers[0][29] ,
         \registers[0][28] , \registers[0][27] , \registers[0][26] ,
         \registers[0][25] , \registers[0][24] , \registers[0][23] ,
         \registers[0][22] , \registers[0][21] , \registers[0][20] ,
         \registers[0][19] , \registers[0][18] , \registers[0][17] ,
         \registers[0][16] , \registers[0][15] , \registers[0][14] ,
         \registers[0][13] , \registers[0][12] , \registers[0][11] ,
         \registers[0][10] , \registers[0][9] , \registers[0][8] ,
         \registers[0][7] , \registers[0][6] , \registers[0][5] ,
         \registers[0][4] , \registers[0][3] , \registers[0][2] ,
         \registers[0][1] , \registers[0][0] , \registers[1][31] ,
         \registers[1][30] , \registers[1][29] , \registers[1][28] ,
         \registers[1][27] , \registers[1][26] , \registers[1][25] ,
         \registers[1][24] , \registers[1][23] , \registers[1][22] ,
         \registers[1][21] , \registers[1][20] , \registers[1][19] ,
         \registers[1][18] , \registers[1][17] , \registers[1][16] ,
         \registers[1][15] , \registers[1][14] , \registers[1][13] ,
         \registers[1][12] , \registers[1][11] , \registers[1][10] ,
         \registers[1][9] , \registers[1][8] , \registers[1][7] ,
         \registers[1][6] , \registers[1][5] , \registers[1][4] ,
         \registers[1][3] , \registers[1][2] , \registers[1][1] ,
         \registers[1][0] , \registers[2][31] , \registers[2][30] ,
         \registers[2][29] , \registers[2][28] , \registers[2][27] ,
         \registers[2][26] , \registers[2][25] , \registers[2][24] ,
         \registers[2][23] , \registers[2][22] , \registers[2][21] ,
         \registers[2][20] , \registers[2][19] , \registers[2][18] ,
         \registers[2][17] , \registers[2][16] , \registers[2][15] ,
         \registers[2][14] , \registers[2][13] , \registers[2][12] ,
         \registers[2][11] , \registers[2][10] , \registers[2][9] ,
         \registers[2][8] , \registers[2][7] , \registers[2][6] ,
         \registers[2][5] , \registers[2][4] , \registers[2][3] ,
         \registers[2][2] , \registers[2][1] , \registers[2][0] ,
         \registers[3][31] , \registers[3][30] , \registers[3][29] ,
         \registers[3][28] , \registers[3][27] , \registers[3][26] ,
         \registers[3][25] , \registers[3][24] , \registers[3][23] ,
         \registers[3][22] , \registers[3][21] , \registers[3][20] ,
         \registers[3][19] , \registers[3][18] , \registers[3][17] ,
         \registers[3][16] , \registers[3][15] , \registers[3][14] ,
         \registers[3][13] , \registers[3][12] , \registers[3][11] ,
         \registers[3][10] , \registers[3][9] , \registers[3][8] ,
         \registers[3][7] , \registers[3][6] , \registers[3][5] ,
         \registers[3][4] , \registers[3][3] , \registers[3][2] ,
         \registers[3][1] , \registers[3][0] , \registers[4][31] ,
         \registers[4][30] , \registers[4][29] , \registers[4][28] ,
         \registers[4][27] , \registers[4][26] , \registers[4][25] ,
         \registers[4][24] , \registers[4][23] , \registers[4][22] ,
         \registers[4][21] , \registers[4][20] , \registers[4][19] ,
         \registers[4][18] , \registers[4][17] , \registers[4][16] ,
         \registers[4][15] , \registers[4][14] , \registers[4][13] ,
         \registers[4][12] , \registers[4][11] , \registers[4][10] ,
         \registers[4][9] , \registers[4][8] , \registers[4][7] ,
         \registers[4][6] , \registers[4][5] , \registers[4][4] ,
         \registers[4][3] , \registers[4][2] , \registers[4][1] ,
         \registers[4][0] , \registers[5][31] , \registers[5][30] ,
         \registers[5][29] , \registers[5][28] , \registers[5][27] ,
         \registers[5][26] , \registers[5][25] , \registers[5][24] ,
         \registers[5][23] , \registers[5][22] , \registers[5][21] ,
         \registers[5][20] , \registers[5][19] , \registers[5][18] ,
         \registers[5][17] , \registers[5][16] , \registers[5][15] ,
         \registers[5][14] , \registers[5][13] , \registers[5][12] ,
         \registers[5][11] , \registers[5][10] , \registers[5][9] ,
         \registers[5][8] , \registers[5][7] , \registers[5][6] ,
         \registers[5][5] , \registers[5][4] , \registers[5][3] ,
         \registers[5][2] , \registers[5][1] , \registers[5][0] ,
         \registers[6][31] , \registers[6][30] , \registers[6][29] ,
         \registers[6][28] , \registers[6][27] , \registers[6][26] ,
         \registers[6][25] , \registers[6][24] , \registers[6][23] ,
         \registers[6][22] , \registers[6][21] , \registers[6][20] ,
         \registers[6][19] , \registers[6][18] , \registers[6][17] ,
         \registers[6][16] , \registers[6][15] , \registers[6][14] ,
         \registers[6][13] , \registers[6][12] , \registers[6][11] ,
         \registers[6][10] , \registers[6][9] , \registers[6][8] ,
         \registers[6][7] , \registers[6][6] , \registers[6][5] ,
         \registers[6][4] , \registers[6][3] , \registers[6][2] ,
         \registers[6][1] , \registers[6][0] , \registers[7][31] ,
         \registers[7][30] , \registers[7][29] , \registers[7][28] ,
         \registers[7][27] , \registers[7][26] , \registers[7][25] ,
         \registers[7][24] , \registers[7][23] , \registers[7][22] ,
         \registers[7][21] , \registers[7][20] , \registers[7][19] ,
         \registers[7][18] , \registers[7][17] , \registers[7][16] ,
         \registers[7][15] , \registers[7][14] , \registers[7][13] ,
         \registers[7][12] , \registers[7][11] , \registers[7][10] ,
         \registers[7][9] , \registers[7][8] , \registers[7][7] ,
         \registers[7][6] , \registers[7][5] , \registers[7][4] ,
         \registers[7][3] , \registers[7][2] , \registers[7][1] ,
         \registers[7][0] , \registers[8][31] , \registers[8][30] ,
         \registers[8][29] , \registers[8][28] , \registers[8][27] ,
         \registers[8][26] , \registers[8][25] , \registers[8][24] ,
         \registers[8][23] , \registers[8][22] , \registers[8][21] ,
         \registers[8][20] , \registers[8][19] , \registers[8][18] ,
         \registers[8][17] , \registers[8][16] , \registers[8][15] ,
         \registers[8][14] , \registers[8][13] , \registers[8][12] ,
         \registers[8][11] , \registers[8][10] , \registers[8][9] ,
         \registers[8][8] , \registers[8][7] , \registers[8][6] ,
         \registers[8][5] , \registers[8][4] , \registers[8][3] ,
         \registers[8][2] , \registers[8][1] , \registers[8][0] ,
         \registers[9][31] , \registers[9][30] , \registers[9][29] ,
         \registers[9][28] , \registers[9][27] , \registers[9][26] ,
         \registers[9][25] , \registers[9][24] , \registers[9][23] ,
         \registers[9][22] , \registers[9][21] , \registers[9][20] ,
         \registers[9][19] , \registers[9][18] , \registers[9][17] ,
         \registers[9][16] , \registers[9][15] , \registers[9][14] ,
         \registers[9][13] , \registers[9][12] , \registers[9][11] ,
         \registers[9][10] , \registers[9][9] , \registers[9][8] ,
         \registers[9][7] , \registers[9][6] , \registers[9][5] ,
         \registers[9][4] , \registers[9][3] , \registers[9][2] ,
         \registers[9][1] , \registers[9][0] , \registers[10][31] ,
         \registers[10][30] , \registers[10][29] , \registers[10][28] ,
         \registers[10][27] , \registers[10][26] , \registers[10][25] ,
         \registers[10][24] , \registers[10][23] , \registers[10][22] ,
         \registers[10][21] , \registers[10][20] , \registers[10][19] ,
         \registers[10][18] , \registers[10][17] , \registers[10][16] ,
         \registers[10][15] , \registers[10][14] , \registers[10][13] ,
         \registers[10][12] , \registers[10][11] , \registers[10][10] ,
         \registers[10][9] , \registers[10][8] , \registers[10][7] ,
         \registers[10][6] , \registers[10][5] , \registers[10][4] ,
         \registers[10][3] , \registers[10][2] , \registers[10][1] ,
         \registers[10][0] , \registers[11][31] , \registers[11][30] ,
         \registers[11][29] , \registers[11][28] , \registers[11][27] ,
         \registers[11][26] , \registers[11][25] , \registers[11][24] ,
         \registers[11][23] , \registers[11][22] , \registers[11][21] ,
         \registers[11][20] , \registers[11][19] , \registers[11][18] ,
         \registers[11][17] , \registers[11][16] , \registers[11][15] ,
         \registers[11][14] , \registers[11][13] , \registers[11][12] ,
         \registers[11][11] , \registers[11][10] , \registers[11][9] ,
         \registers[11][8] , \registers[11][7] , \registers[11][6] ,
         \registers[11][5] , \registers[11][4] , \registers[11][3] ,
         \registers[11][2] , \registers[11][1] , \registers[11][0] ,
         \registers[12][31] , \registers[12][30] , \registers[12][29] ,
         \registers[12][28] , \registers[12][27] , \registers[12][26] ,
         \registers[12][25] , \registers[12][24] , \registers[12][23] ,
         \registers[12][22] , \registers[12][21] , \registers[12][20] ,
         \registers[12][19] , \registers[12][18] , \registers[12][17] ,
         \registers[12][16] , \registers[12][15] , \registers[12][14] ,
         \registers[12][13] , \registers[12][12] , \registers[12][11] ,
         \registers[12][10] , \registers[12][9] , \registers[12][8] ,
         \registers[12][7] , \registers[12][6] , \registers[12][5] ,
         \registers[12][4] , \registers[12][3] , \registers[12][2] ,
         \registers[12][1] , \registers[12][0] , \registers[13][31] ,
         \registers[13][30] , \registers[13][29] , \registers[13][28] ,
         \registers[13][27] , \registers[13][26] , \registers[13][25] ,
         \registers[13][24] , \registers[13][23] , \registers[13][22] ,
         \registers[13][21] , \registers[13][20] , \registers[13][19] ,
         \registers[13][18] , \registers[13][17] , \registers[13][16] ,
         \registers[13][15] , \registers[13][14] , \registers[13][13] ,
         \registers[13][12] , \registers[13][11] , \registers[13][10] ,
         \registers[13][9] , \registers[13][8] , \registers[13][7] ,
         \registers[13][6] , \registers[13][5] , \registers[13][4] ,
         \registers[13][3] , \registers[13][2] , \registers[13][1] ,
         \registers[13][0] , \registers[14][31] , \registers[14][30] ,
         \registers[14][29] , \registers[14][28] , \registers[14][27] ,
         \registers[14][26] , \registers[14][25] , \registers[14][24] ,
         \registers[14][23] , \registers[14][22] , \registers[14][21] ,
         \registers[14][20] , \registers[14][19] , \registers[14][18] ,
         \registers[14][17] , \registers[14][16] , \registers[14][15] ,
         \registers[14][14] , \registers[14][13] , \registers[14][12] ,
         \registers[14][11] , \registers[14][10] , \registers[14][9] ,
         \registers[14][8] , \registers[14][7] , \registers[14][6] ,
         \registers[14][5] , \registers[14][4] , \registers[14][3] ,
         \registers[14][2] , \registers[14][1] , \registers[14][0] ,
         \registers[15][31] , \registers[15][30] , \registers[15][29] ,
         \registers[15][28] , \registers[15][27] , \registers[15][26] ,
         \registers[15][25] , \registers[15][24] , \registers[15][23] ,
         \registers[15][22] , \registers[15][21] , \registers[15][20] ,
         \registers[15][19] , \registers[15][18] , \registers[15][17] ,
         \registers[15][16] , \registers[15][15] , \registers[15][14] ,
         \registers[15][13] , \registers[15][12] , \registers[15][11] ,
         \registers[15][10] , \registers[15][9] , \registers[15][8] ,
         \registers[15][7] , \registers[15][6] , \registers[15][5] ,
         \registers[15][4] , \registers[15][3] , \registers[15][2] ,
         \registers[15][1] , \registers[15][0] , \registers[16][31] ,
         \registers[16][30] , \registers[16][29] , \registers[16][28] ,
         \registers[16][27] , \registers[16][26] , \registers[16][25] ,
         \registers[16][24] , \registers[16][23] , \registers[16][22] ,
         \registers[16][21] , \registers[16][20] , \registers[16][19] ,
         \registers[16][18] , \registers[16][17] , \registers[16][16] ,
         \registers[16][15] , \registers[16][14] , \registers[16][13] ,
         \registers[16][12] , \registers[16][11] , \registers[16][10] ,
         \registers[16][9] , \registers[16][8] , \registers[16][7] ,
         \registers[16][6] , \registers[16][5] , \registers[16][4] ,
         \registers[16][3] , \registers[16][2] , \registers[16][1] ,
         \registers[16][0] , \registers[17][31] , \registers[17][30] ,
         \registers[17][29] , \registers[17][28] , \registers[17][27] ,
         \registers[17][26] , \registers[17][25] , \registers[17][24] ,
         \registers[17][23] , \registers[17][22] , \registers[17][21] ,
         \registers[17][20] , \registers[17][19] , \registers[17][18] ,
         \registers[17][17] , \registers[17][16] , \registers[17][15] ,
         \registers[17][14] , \registers[17][13] , \registers[17][12] ,
         \registers[17][11] , \registers[17][10] , \registers[17][9] ,
         \registers[17][8] , \registers[17][7] , \registers[17][6] ,
         \registers[17][5] , \registers[17][4] , \registers[17][3] ,
         \registers[17][2] , \registers[17][1] , \registers[17][0] ,
         \registers[18][31] , \registers[18][30] , \registers[18][29] ,
         \registers[18][28] , \registers[18][27] , \registers[18][26] ,
         \registers[18][25] , \registers[18][24] , \registers[18][23] ,
         \registers[18][22] , \registers[18][21] , \registers[18][20] ,
         \registers[18][19] , \registers[18][18] , \registers[18][17] ,
         \registers[18][16] , \registers[18][15] , \registers[18][14] ,
         \registers[18][13] , \registers[18][12] , \registers[18][11] ,
         \registers[18][10] , \registers[18][9] , \registers[18][8] ,
         \registers[18][7] , \registers[18][6] , \registers[18][5] ,
         \registers[18][4] , \registers[18][3] , \registers[18][2] ,
         \registers[18][1] , \registers[18][0] , \registers[19][31] ,
         \registers[19][30] , \registers[19][29] , \registers[19][28] ,
         \registers[19][27] , \registers[19][26] , \registers[19][25] ,
         \registers[19][24] , \registers[19][23] , \registers[19][22] ,
         \registers[19][21] , \registers[19][20] , \registers[19][19] ,
         \registers[19][18] , \registers[19][17] , \registers[19][16] ,
         \registers[19][15] , \registers[19][14] , \registers[19][13] ,
         \registers[19][12] , \registers[19][11] , \registers[19][10] ,
         \registers[19][9] , \registers[19][8] , \registers[19][7] ,
         \registers[19][6] , \registers[19][5] , \registers[19][4] ,
         \registers[19][3] , \registers[19][2] , \registers[19][1] ,
         \registers[19][0] , \registers[20][31] , \registers[20][30] ,
         \registers[20][29] , \registers[20][28] , \registers[20][27] ,
         \registers[20][26] , \registers[20][25] , \registers[20][24] ,
         \registers[20][23] , \registers[20][22] , \registers[20][21] ,
         \registers[20][20] , \registers[20][19] , \registers[20][18] ,
         \registers[20][17] , \registers[20][16] , \registers[20][15] ,
         \registers[20][14] , \registers[20][13] , \registers[20][12] ,
         \registers[20][11] , \registers[20][10] , \registers[20][9] ,
         \registers[20][8] , \registers[20][7] , \registers[20][6] ,
         \registers[20][5] , \registers[20][4] , \registers[20][3] ,
         \registers[20][2] , \registers[20][1] , \registers[20][0] ,
         \registers[21][31] , \registers[21][30] , \registers[21][29] ,
         \registers[21][28] , \registers[21][27] , \registers[21][26] ,
         \registers[21][25] , \registers[21][24] , \registers[21][23] ,
         \registers[21][22] , \registers[21][21] , \registers[21][20] ,
         \registers[21][19] , \registers[21][18] , \registers[21][17] ,
         \registers[21][16] , \registers[21][15] , \registers[21][14] ,
         \registers[21][13] , \registers[21][12] , \registers[21][11] ,
         \registers[21][10] , \registers[21][9] , \registers[21][8] ,
         \registers[21][7] , \registers[21][6] , \registers[21][5] ,
         \registers[21][4] , \registers[21][3] , \registers[21][2] ,
         \registers[21][1] , \registers[21][0] , \registers[22][31] ,
         \registers[22][30] , \registers[22][29] , \registers[22][28] ,
         \registers[22][27] , \registers[22][26] , \registers[22][25] ,
         \registers[22][24] , \registers[22][23] , \registers[22][22] ,
         \registers[22][21] , \registers[22][20] , \registers[22][19] ,
         \registers[22][18] , \registers[22][17] , \registers[22][16] ,
         \registers[22][15] , \registers[22][14] , \registers[22][13] ,
         \registers[22][12] , \registers[22][11] , \registers[22][10] ,
         \registers[22][9] , \registers[22][8] , \registers[22][7] ,
         \registers[22][6] , \registers[22][5] , \registers[22][4] ,
         \registers[22][3] , \registers[22][2] , \registers[22][1] ,
         \registers[22][0] , \registers[23][31] , \registers[23][30] ,
         \registers[23][29] , \registers[23][28] , \registers[23][27] ,
         \registers[23][26] , \registers[23][25] , \registers[23][24] ,
         \registers[23][23] , \registers[23][22] , \registers[23][21] ,
         \registers[23][20] , \registers[23][19] , \registers[23][18] ,
         \registers[23][17] , \registers[23][16] , \registers[23][15] ,
         \registers[23][14] , \registers[23][13] , \registers[23][12] ,
         \registers[23][11] , \registers[23][10] , \registers[23][9] ,
         \registers[23][8] , \registers[23][7] , \registers[23][6] ,
         \registers[23][5] , \registers[23][4] , \registers[23][3] ,
         \registers[23][2] , \registers[23][1] , \registers[23][0] ,
         \registers[24][31] , \registers[24][30] , \registers[24][29] ,
         \registers[24][28] , \registers[24][27] , \registers[24][26] ,
         \registers[24][25] , \registers[24][24] , \registers[24][23] ,
         \registers[24][22] , \registers[24][21] , \registers[24][20] ,
         \registers[24][19] , \registers[24][18] , \registers[24][17] ,
         \registers[24][16] , \registers[24][15] , \registers[24][14] ,
         \registers[24][13] , \registers[24][12] , \registers[24][11] ,
         \registers[24][10] , \registers[24][9] , \registers[24][8] ,
         \registers[24][7] , \registers[24][6] , \registers[24][5] ,
         \registers[24][4] , \registers[24][3] , \registers[24][2] ,
         \registers[24][1] , \registers[24][0] , \registers[25][31] ,
         \registers[25][30] , \registers[25][29] , \registers[25][28] ,
         \registers[25][27] , \registers[25][26] , \registers[25][25] ,
         \registers[25][24] , \registers[25][23] , \registers[25][22] ,
         \registers[25][21] , \registers[25][20] , \registers[25][19] ,
         \registers[25][18] , \registers[25][17] , \registers[25][16] ,
         \registers[25][15] , \registers[25][14] , \registers[25][13] ,
         \registers[25][12] , \registers[25][11] , \registers[25][10] ,
         \registers[25][9] , \registers[25][8] , \registers[25][7] ,
         \registers[25][6] , \registers[25][5] , \registers[25][4] ,
         \registers[25][3] , \registers[25][2] , \registers[25][1] ,
         \registers[25][0] , \registers[26][31] , \registers[26][30] ,
         \registers[26][29] , \registers[26][28] , \registers[26][27] ,
         \registers[26][26] , \registers[26][25] , \registers[26][24] ,
         \registers[26][23] , \registers[26][22] , \registers[26][21] ,
         \registers[26][20] , \registers[26][19] , \registers[26][18] ,
         \registers[26][17] , \registers[26][16] , \registers[26][15] ,
         \registers[26][14] , \registers[26][13] , \registers[26][12] ,
         \registers[26][11] , \registers[26][10] , \registers[26][9] ,
         \registers[26][8] , \registers[26][7] , \registers[26][6] ,
         \registers[26][5] , \registers[26][4] , \registers[26][3] ,
         \registers[26][2] , \registers[26][1] , \registers[26][0] ,
         \registers[27][31] , \registers[27][30] , \registers[27][29] ,
         \registers[27][28] , \registers[27][27] , \registers[27][26] ,
         \registers[27][25] , \registers[27][24] , \registers[27][23] ,
         \registers[27][22] , \registers[27][21] , \registers[27][20] ,
         \registers[27][19] , \registers[27][18] , \registers[27][17] ,
         \registers[27][16] , \registers[27][15] , \registers[27][14] ,
         \registers[27][13] , \registers[27][12] , \registers[27][11] ,
         \registers[27][10] , \registers[27][9] , \registers[27][8] ,
         \registers[27][7] , \registers[27][6] , \registers[27][5] ,
         \registers[27][4] , \registers[27][3] , \registers[27][2] ,
         \registers[27][1] , \registers[27][0] , \registers[28][31] ,
         \registers[28][30] , \registers[28][29] , \registers[28][28] ,
         \registers[28][27] , \registers[28][26] , \registers[28][25] ,
         \registers[28][24] , \registers[28][23] , \registers[28][22] ,
         \registers[28][21] , \registers[28][20] , \registers[28][19] ,
         \registers[28][18] , \registers[28][17] , \registers[28][16] ,
         \registers[28][15] , \registers[28][14] , \registers[28][13] ,
         \registers[28][12] , \registers[28][11] , \registers[28][10] ,
         \registers[28][9] , \registers[28][8] , \registers[28][7] ,
         \registers[28][6] , \registers[28][5] , \registers[28][4] ,
         \registers[28][3] , \registers[28][2] , \registers[28][1] ,
         \registers[28][0] , \registers[29][31] , \registers[29][30] ,
         \registers[29][29] , \registers[29][28] , \registers[29][27] ,
         \registers[29][26] , \registers[29][25] , \registers[29][24] ,
         \registers[29][23] , \registers[29][22] , \registers[29][21] ,
         \registers[29][20] , \registers[29][19] , \registers[29][18] ,
         \registers[29][17] , \registers[29][16] , \registers[29][15] ,
         \registers[29][14] , \registers[29][13] , \registers[29][12] ,
         \registers[29][11] , \registers[29][10] , \registers[29][9] ,
         \registers[29][8] , \registers[29][7] , \registers[29][6] ,
         \registers[29][5] , \registers[29][4] , \registers[29][3] ,
         \registers[29][2] , \registers[29][1] , \registers[29][0] ,
         \registers[30][31] , \registers[30][30] , \registers[30][29] ,
         \registers[30][28] , \registers[30][27] , \registers[30][26] ,
         \registers[30][25] , \registers[30][24] , \registers[30][23] ,
         \registers[30][22] , \registers[30][21] , \registers[30][20] ,
         \registers[30][19] , \registers[30][18] , \registers[30][17] ,
         \registers[30][16] , \registers[30][15] , \registers[30][14] ,
         \registers[30][13] , \registers[30][12] , \registers[30][11] ,
         \registers[30][10] , \registers[30][9] , \registers[30][8] ,
         \registers[30][7] , \registers[30][6] , \registers[30][5] ,
         \registers[30][4] , \registers[30][3] , \registers[30][2] ,
         \registers[30][1] , \registers[30][0] , \registers[31][31] ,
         \registers[31][30] , \registers[31][29] , \registers[31][28] ,
         \registers[31][27] , \registers[31][26] , \registers[31][25] ,
         \registers[31][24] , \registers[31][23] , \registers[31][22] ,
         \registers[31][21] , \registers[31][20] , \registers[31][19] ,
         \registers[31][18] , \registers[31][17] , \registers[31][16] ,
         \registers[31][15] , \registers[31][14] , \registers[31][13] ,
         \registers[31][12] , \registers[31][11] , \registers[31][10] ,
         \registers[31][9] , \registers[31][8] , \registers[31][7] ,
         \registers[31][6] , \registers[31][5] , \registers[31][4] ,
         \registers[31][3] , \registers[31][2] , \registers[31][1] ,
         \registers[31][0] , n2956, n2958, n2960, n2962, n2964, n2966, n2968,
         n2970, n2972, n2974, n2976, n2978, n2980, n2982, n2984, n2986, n2988,
         n2990, n2992, n2994, n2996, n2998, n3000, n3002, n3004, n3006, n3008,
         n3010, n3012, n3014, n3016, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n675, n1684, n1685, n1688, n1690,
         n1692, n1694, n1696, n1698, n1700, n1702, n1704, n1706, n1708, n1710,
         n1712, n1714, n1716, n1718, n1720, n1722, n1724, n1726, n1728, n1730,
         n1732, n1734, n1736, n1738, n1740, n1742, n1744, n1746, n1748, n1750,
         n1751, n1786, n1787, n1788, n1821, n1822, n1823, n1856, n1857, n1858,
         n1859, n1860, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n2031, n2032, n2066,
         n2100, n2582, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2755, n2756,
         n2757, n2790, n2824, n2825, n2858, n2859, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2957,
         n2959, n2961, n2963, n2965, n2967, n2969, n2973, n2975, n2977, n2979,
         n2981, n2983, n2985, n2987, n2989, n2991, n2993, n2995, n2997, n2999,
         n3001, n3003, n3005, n3007, n3009, n3011, n3013, n3015, n3017, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4182, n4183, n4184, n4217, n4251, n4252, n4285, n4286, n4319, n4320,
         n4321, n4354, n4355, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2583, n2618, n2652, n2686,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2860,
         n2895, n2929, n2971, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4356, n4390, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872;

  DFFR_X1 \registers_reg[0][31]  ( .D(n4138), .CK(n675), .RN(n6836), .Q(
        \registers[0][31] ), .QN(n5763) );
  DFFR_X1 \registers_reg[0][30]  ( .D(n4137), .CK(n675), .RN(n6831), .Q(
        \registers[0][30] ), .QN(n5762) );
  DFFR_X1 \registers_reg[0][29]  ( .D(n4136), .CK(n675), .RN(n6825), .Q(
        \registers[0][29] ), .QN(n5783) );
  DFFR_X1 \registers_reg[0][28]  ( .D(n4135), .CK(n675), .RN(n6820), .Q(
        \registers[0][28] ), .QN(n4295) );
  DFFR_X1 \registers_reg[0][27]  ( .D(n4134), .CK(n675), .RN(n6839), .Q(
        \registers[0][27] ), .QN(n5761) );
  DFFR_X1 \registers_reg[0][26]  ( .D(n4133), .CK(n675), .RN(n6811), .Q(
        \registers[0][26] ), .QN(n5782) );
  DFFR_X1 \registers_reg[0][25]  ( .D(n4132), .CK(n675), .RN(n6814), .Q(
        \registers[0][25] ), .QN(n5760) );
  DFFR_X1 \registers_reg[0][24]  ( .D(n4131), .CK(n675), .RN(n6806), .Q(
        \registers[0][24] ), .QN(n5759) );
  DFFR_X1 \registers_reg[0][23]  ( .D(n4130), .CK(n675), .RN(n6842), .Q(
        \registers[0][23] ), .QN(n5781) );
  DFFR_X1 \registers_reg[0][22]  ( .D(n4129), .CK(n675), .RN(n6795), .Q(
        \registers[0][22] ), .QN(n4390) );
  DFFR_X1 \registers_reg[0][21]  ( .D(n4128), .CK(n675), .RN(n6798), .Q(
        \registers[0][21] ), .QN(n4294) );
  DFFR_X1 \registers_reg[0][20]  ( .D(n4127), .CK(n675), .RN(n6789), .Q(
        \registers[0][20] ), .QN(n5780) );
  DFFR_X1 \registers_reg[0][19]  ( .D(n4126), .CK(n675), .RN(n6845), .Q(
        \registers[0][19] ), .QN(n4293) );
  DFFR_X1 \registers_reg[0][18]  ( .D(n4125), .CK(n675), .RN(n6778), .Q(
        \registers[0][18] ), .QN(n4292) );
  DFFR_X1 \registers_reg[0][17]  ( .D(n4124), .CK(n675), .RN(n6781), .Q(
        \registers[0][17] ), .QN(n5779) );
  DFFR_X1 \registers_reg[0][16]  ( .D(n4123), .CK(n675), .RN(n6772), .Q(
        \registers[0][16] ), .QN(n4356) );
  DFFR_X1 \registers_reg[0][15]  ( .D(n4122), .CK(n675), .RN(n6848), .Q(
        \registers[0][15] ), .QN(n4353) );
  DFFR_X1 \registers_reg[0][14]  ( .D(n4121), .CK(n675), .RN(n6828), .Q(
        \registers[0][14] ), .QN(n5778) );
  DFFR_X1 \registers_reg[0][13]  ( .D(n4120), .CK(n675), .RN(n6822), .Q(
        \registers[0][13] ), .QN(n4352) );
  DFFR_X1 \registers_reg[0][12]  ( .D(n4119), .CK(n675), .RN(n6817), .Q(
        \registers[0][12] ), .QN(n4351) );
  DFFR_X1 \registers_reg[0][11]  ( .D(n4118), .CK(n675), .RN(n6850), .Q(
        \registers[0][11] ), .QN(n5777) );
  DFFR_X1 \registers_reg[0][10]  ( .D(n4117), .CK(n675), .RN(n6809), .Q(
        \registers[0][10] ), .QN(n4291) );
  DFFR_X1 \registers_reg[0][9]  ( .D(n4116), .CK(n675), .RN(n6800), .Q(
        \registers[0][9] ), .QN(n4350) );
  DFFR_X1 \registers_reg[0][8]  ( .D(n4115), .CK(n675), .RN(n6803), .Q(
        \registers[0][8] ), .QN(n5776) );
  DFFR_X1 \registers_reg[0][7]  ( .D(n4114), .CK(n675), .RN(n6853), .Q(
        \registers[0][7] ), .QN(n4349) );
  DFFR_X1 \registers_reg[0][6]  ( .D(n4113), .CK(n675), .RN(n6792), .Q(
        \registers[0][6] ), .QN(n4348) );
  DFFR_X1 \registers_reg[0][5]  ( .D(n4112), .CK(n675), .RN(n6784), .Q(
        \registers[0][5] ), .QN(n5775) );
  DFFR_X1 \registers_reg[0][4]  ( .D(n4111), .CK(n675), .RN(n6786), .Q(
        \registers[0][4] ), .QN(n4347) );
  DFFR_X1 \registers_reg[0][3]  ( .D(n4110), .CK(n675), .RN(n6834), .Q(
        \registers[0][3] ), .QN(n4290) );
  DFFR_X1 \registers_reg[0][2]  ( .D(n4109), .CK(n675), .RN(n6775), .Q(
        \registers[0][2] ), .QN(n5774) );
  DFFR_X1 \registers_reg[0][1]  ( .D(n4108), .CK(n675), .RN(n6770), .Q(
        \registers[0][1] ), .QN(n4289) );
  DFFR_X1 \registers_reg[0][0]  ( .D(n4107), .CK(n675), .RN(n6856), .Q(
        \registers[0][0] ), .QN(n4288) );
  DFFR_X1 \registers_reg[1][31]  ( .D(n4106), .CK(n675), .RN(n6836), .Q(
        \registers[1][31] ), .QN(n2770) );
  DFFR_X1 \registers_reg[1][30]  ( .D(n4105), .CK(n675), .RN(n6831), .Q(
        \registers[1][30] ), .QN(n2769) );
  DFFR_X1 \registers_reg[1][29]  ( .D(n4104), .CK(n675), .RN(n6825), .Q(
        \registers[1][29] ), .QN(n2791) );
  DFFR_X1 \registers_reg[1][28]  ( .D(n4103), .CK(n675), .RN(n6820), .Q(
        \registers[1][28] ), .QN(n2568) );
  DFFR_X1 \registers_reg[1][27]  ( .D(n4102), .CK(n675), .RN(n6839), .Q(
        \registers[1][27] ), .QN(n2768) );
  DFFR_X1 \registers_reg[1][26]  ( .D(n4101), .CK(n675), .RN(n6811), .Q(
        \registers[1][26] ), .QN(n2789) );
  DFFR_X1 \registers_reg[1][25]  ( .D(n4100), .CK(n675), .RN(n6814), .Q(
        \registers[1][25] ), .QN(n2767) );
  DFFR_X1 \registers_reg[1][24]  ( .D(n4099), .CK(n675), .RN(n6806), .Q(
        \registers[1][24] ), .QN(n2766) );
  DFFR_X1 \registers_reg[1][23]  ( .D(n4098), .CK(n675), .RN(n6842), .Q(
        \registers[1][23] ), .QN(n2788) );
  DFFR_X1 \registers_reg[1][22]  ( .D(n4097), .CK(n675), .RN(n6795), .Q(
        \registers[1][22] ), .QN(n2765) );
  DFFR_X1 \registers_reg[1][21]  ( .D(n4096), .CK(n675), .RN(n6797), .Q(
        \registers[1][21] ), .QN(n2567) );
  DFFR_X1 \registers_reg[1][20]  ( .D(n4095), .CK(n675), .RN(n6789), .Q(
        \registers[1][20] ), .QN(n2787) );
  DFFR_X1 \registers_reg[1][19]  ( .D(n4094), .CK(n675), .RN(n6845), .Q(
        \registers[1][19] ), .QN(n2566) );
  DFFR_X1 \registers_reg[1][18]  ( .D(n4093), .CK(n675), .RN(n6778), .Q(
        \registers[1][18] ), .QN(n2565) );
  DFFR_X1 \registers_reg[1][17]  ( .D(n4092), .CK(n675), .RN(n6781), .Q(
        \registers[1][17] ), .QN(n2786) );
  DFFR_X1 \registers_reg[1][16]  ( .D(n4091), .CK(n675), .RN(n6772), .Q(
        \registers[1][16] ), .QN(n2764) );
  DFFR_X1 \registers_reg[1][15]  ( .D(n4090), .CK(n675), .RN(n6848), .Q(
        \registers[1][15] ), .QN(n2763) );
  DFFR_X1 \registers_reg[1][14]  ( .D(n4089), .CK(n675), .RN(n6828), .Q(
        \registers[1][14] ), .QN(n2785) );
  DFFR_X1 \registers_reg[1][13]  ( .D(n4088), .CK(n675), .RN(n6822), .Q(
        \registers[1][13] ), .QN(n2762) );
  DFFR_X1 \registers_reg[1][12]  ( .D(n4087), .CK(n675), .RN(n6817), .Q(
        \registers[1][12] ), .QN(n2761) );
  DFFR_X1 \registers_reg[1][11]  ( .D(n4086), .CK(n675), .RN(n6850), .Q(
        \registers[1][11] ), .QN(n2784) );
  DFFR_X1 \registers_reg[1][10]  ( .D(n4085), .CK(n675), .RN(n6809), .Q(
        \registers[1][10] ), .QN(n2564) );
  DFFR_X1 \registers_reg[1][9]  ( .D(n4084), .CK(n675), .RN(n6800), .Q(
        \registers[1][9] ), .QN(n2760) );
  DFFR_X1 \registers_reg[1][8]  ( .D(n4083), .CK(n675), .RN(n6803), .Q(
        \registers[1][8] ), .QN(n2783) );
  DFFR_X1 \registers_reg[1][7]  ( .D(n4082), .CK(n675), .RN(n6853), .Q(
        \registers[1][7] ), .QN(n2759) );
  DFFR_X1 \registers_reg[1][6]  ( .D(n4081), .CK(n675), .RN(n6792), .Q(
        \registers[1][6] ), .QN(n2758) );
  DFFR_X1 \registers_reg[1][5]  ( .D(n4080), .CK(n675), .RN(n6784), .Q(
        \registers[1][5] ), .QN(n2782) );
  DFFR_X1 \registers_reg[1][4]  ( .D(n4079), .CK(n675), .RN(n6786), .Q(
        \registers[1][4] ), .QN(n2754) );
  DFFR_X1 \registers_reg[1][3]  ( .D(n4078), .CK(n675), .RN(n6833), .Q(
        \registers[1][3] ), .QN(n2563) );
  DFFR_X1 \registers_reg[1][2]  ( .D(n4077), .CK(n675), .RN(n6775), .Q(
        \registers[1][2] ), .QN(n2781) );
  DFFR_X1 \registers_reg[1][1]  ( .D(n4076), .CK(n675), .RN(n6770), .Q(
        \registers[1][1] ), .QN(n2562) );
  DFFR_X1 \registers_reg[1][0]  ( .D(n4075), .CK(n675), .RN(n6856), .Q(
        \registers[1][0] ), .QN(n2561) );
  DFFR_X1 \registers_reg[2][31]  ( .D(n4074), .CK(n675), .RN(n6836), .Q(
        \registers[2][31] ), .QN(n2731) );
  DFFR_X1 \registers_reg[2][30]  ( .D(n4073), .CK(n675), .RN(n6831), .Q(
        \registers[2][30] ), .QN(n2730) );
  DFFR_X1 \registers_reg[2][29]  ( .D(n4072), .CK(n675), .RN(n6825), .Q(
        \registers[2][29] ), .QN(n2729) );
  DFFR_X1 \registers_reg[2][28]  ( .D(n4071), .CK(n675), .RN(n6820), .Q(
        \registers[2][28] ), .QN(n2728) );
  DFFR_X1 \registers_reg[2][27]  ( .D(n4070), .CK(n675), .RN(n6839), .Q(
        \registers[2][27] ), .QN(n4212) );
  DFFR_X1 \registers_reg[2][26]  ( .D(n4069), .CK(n675), .RN(n6811), .Q(
        \registers[2][26] ), .QN(n4210) );
  DFFR_X1 \registers_reg[2][25]  ( .D(n4068), .CK(n675), .RN(n6814), .Q(
        \registers[2][25] ), .QN(n4208) );
  DFFR_X1 \registers_reg[2][24]  ( .D(n4067), .CK(n675), .RN(n6806), .Q(
        \registers[2][24] ), .QN(n4206) );
  DFFR_X1 \registers_reg[2][23]  ( .D(n4066), .CK(n675), .RN(n6842), .Q(
        \registers[2][23] ), .QN(n4204) );
  DFFR_X1 \registers_reg[2][22]  ( .D(n4065), .CK(n675), .RN(n6795), .Q(
        \registers[2][22] ), .QN(n4202) );
  DFFR_X1 \registers_reg[2][21]  ( .D(n4064), .CK(n675), .RN(n6797), .Q(
        \registers[2][21] ), .QN(n2727) );
  DFFR_X1 \registers_reg[2][20]  ( .D(n4063), .CK(n675), .RN(n6789), .Q(
        \registers[2][20] ), .QN(n2726) );
  DFFR_X1 \registers_reg[2][19]  ( .D(n4062), .CK(n675), .RN(n6845), .Q(
        \registers[2][19] ), .QN(n2725) );
  DFFR_X1 \registers_reg[2][18]  ( .D(n4061), .CK(n675), .RN(n6778), .Q(
        \registers[2][18] ), .QN(n2724) );
  DFFR_X1 \registers_reg[2][17]  ( .D(n4060), .CK(n675), .RN(n6781), .Q(
        \registers[2][17] ), .QN(n2723) );
  DFFR_X1 \registers_reg[2][16]  ( .D(n4059), .CK(n675), .RN(n6772), .Q(
        \registers[2][16] ), .QN(n2686) );
  DFFR_X1 \registers_reg[2][15]  ( .D(n4058), .CK(n675), .RN(n6847), .Q(
        \registers[2][15] ), .QN(n2652) );
  DFFR_X1 \registers_reg[2][14]  ( .D(n4057), .CK(n675), .RN(n6828), .Q(
        \registers[2][14] ), .QN(n2618) );
  DFFR_X1 \registers_reg[2][13]  ( .D(n4056), .CK(n675), .RN(n6822), .Q(
        \registers[2][13] ), .QN(n2583) );
  DFFR_X1 \registers_reg[2][12]  ( .D(n4055), .CK(n675), .RN(n6817), .Q(
        \registers[2][12] ), .QN(n2581) );
  DFFR_X1 \registers_reg[2][11]  ( .D(n4054), .CK(n675), .RN(n6850), .Q(
        \registers[2][11] ), .QN(n2580) );
  DFFR_X1 \registers_reg[2][10]  ( .D(n4053), .CK(n675), .RN(n6808), .Q(
        \registers[2][10] ), .QN(n2579) );
  DFFR_X1 \registers_reg[2][9]  ( .D(n4052), .CK(n675), .RN(n6800), .Q(
        \registers[2][9] ), .QN(n2578) );
  DFFR_X1 \registers_reg[2][8]  ( .D(n4051), .CK(n675), .RN(n6803), .Q(
        \registers[2][8] ), .QN(n2577) );
  DFFR_X1 \registers_reg[2][7]  ( .D(n4050), .CK(n675), .RN(n6853), .Q(
        \registers[2][7] ), .QN(n2576) );
  DFFR_X1 \registers_reg[2][6]  ( .D(n4049), .CK(n675), .RN(n6792), .Q(
        \registers[2][6] ), .QN(n2575) );
  DFFR_X1 \registers_reg[2][5]  ( .D(n4048), .CK(n675), .RN(n6783), .Q(
        \registers[2][5] ), .QN(n2574) );
  DFFR_X1 \registers_reg[2][4]  ( .D(n4047), .CK(n675), .RN(n6786), .Q(
        \registers[2][4] ), .QN(n2573) );
  DFFR_X1 \registers_reg[2][3]  ( .D(n4046), .CK(n675), .RN(n6833), .Q(
        \registers[2][3] ), .QN(n2572) );
  DFFR_X1 \registers_reg[2][2]  ( .D(n4045), .CK(n675), .RN(n6775), .Q(
        \registers[2][2] ), .QN(n2571) );
  DFFR_X1 \registers_reg[2][1]  ( .D(n4044), .CK(n675), .RN(n6770), .Q(
        \registers[2][1] ), .QN(n2570) );
  DFFR_X1 \registers_reg[2][0]  ( .D(n4043), .CK(n675), .RN(n6856), .Q(
        \registers[2][0] ), .QN(n2569) );
  DFFR_X1 \registers_reg[3][31]  ( .D(n4042), .CK(n675), .RN(n6836), .Q(
        \registers[3][31] ), .QN(n4324) );
  DFFR_X1 \registers_reg[3][30]  ( .D(n4041), .CK(n675), .RN(n6830), .Q(
        \registers[3][30] ), .QN(n4323) );
  DFFR_X1 \registers_reg[3][29]  ( .D(n4040), .CK(n675), .RN(n6825), .Q(
        \registers[3][29] ), .QN(n4322) );
  DFFR_X1 \registers_reg[3][28]  ( .D(n4039), .CK(n675), .RN(n6819), .Q(
        \registers[3][28] ), .QN(n4318) );
  DFFR_X1 \registers_reg[3][27]  ( .D(n4038), .CK(n675), .RN(n6839), .Q(
        \registers[3][27] ), .QN(n5911) );
  DFFR_X1 \registers_reg[3][26]  ( .D(n4037), .CK(n675), .RN(n6811), .Q(
        \registers[3][26] ), .QN(n5909) );
  DFFR_X1 \registers_reg[3][25]  ( .D(n4036), .CK(n675), .RN(n6814), .Q(
        \registers[3][25] ), .QN(n5907) );
  DFFR_X1 \registers_reg[3][24]  ( .D(n4035), .CK(n675), .RN(n6806), .Q(
        \registers[3][24] ), .QN(n5905) );
  DFFR_X1 \registers_reg[3][23]  ( .D(n4034), .CK(n675), .RN(n6842), .Q(
        \registers[3][23] ), .QN(n5903) );
  DFFR_X1 \registers_reg[3][22]  ( .D(n4033), .CK(n675), .RN(n6794), .Q(
        \registers[3][22] ), .QN(n5901) );
  DFFR_X1 \registers_reg[3][21]  ( .D(n4032), .CK(n675), .RN(n6797), .Q(
        \registers[3][21] ), .QN(n4317) );
  DFFR_X1 \registers_reg[3][20]  ( .D(n4031), .CK(n675), .RN(n6789), .Q(
        \registers[3][20] ), .QN(n4316) );
  DFFR_X1 \registers_reg[3][19]  ( .D(n4030), .CK(n675), .RN(n6845), .Q(
        \registers[3][19] ), .QN(n4315) );
  DFFR_X1 \registers_reg[3][18]  ( .D(n4029), .CK(n675), .RN(n6778), .Q(
        \registers[3][18] ), .QN(n4314) );
  DFFR_X1 \registers_reg[3][17]  ( .D(n4028), .CK(n675), .RN(n6781), .Q(
        \registers[3][17] ), .QN(n4313) );
  DFFR_X1 \registers_reg[3][16]  ( .D(n4027), .CK(n675), .RN(n6772), .Q(
        \registers[3][16] ), .QN(n4312) );
  DFFR_X1 \registers_reg[3][15]  ( .D(n4026), .CK(n675), .RN(n6847), .Q(
        \registers[3][15] ), .QN(n4311) );
  DFFR_X1 \registers_reg[3][14]  ( .D(n4025), .CK(n675), .RN(n6828), .Q(
        \registers[3][14] ), .QN(n4310) );
  DFFR_X1 \registers_reg[3][13]  ( .D(n4024), .CK(n675), .RN(n6822), .Q(
        \registers[3][13] ), .QN(n4309) );
  DFFR_X1 \registers_reg[3][12]  ( .D(n4023), .CK(n675), .RN(n6817), .Q(
        \registers[3][12] ), .QN(n4308) );
  DFFR_X1 \registers_reg[3][11]  ( .D(n4022), .CK(n675), .RN(n6850), .Q(
        \registers[3][11] ), .QN(n4307) );
  DFFR_X1 \registers_reg[3][10]  ( .D(n4021), .CK(n675), .RN(n6808), .Q(
        \registers[3][10] ), .QN(n4306) );
  DFFR_X1 \registers_reg[3][9]  ( .D(n4020), .CK(n675), .RN(n6800), .Q(
        \registers[3][9] ), .QN(n4305) );
  DFFR_X1 \registers_reg[3][8]  ( .D(n4019), .CK(n675), .RN(n6803), .Q(
        \registers[3][8] ), .QN(n4304) );
  DFFR_X1 \registers_reg[3][7]  ( .D(n4018), .CK(n675), .RN(n6853), .Q(
        \registers[3][7] ), .QN(n4303) );
  DFFR_X1 \registers_reg[3][6]  ( .D(n4017), .CK(n675), .RN(n6792), .Q(
        \registers[3][6] ), .QN(n4302) );
  DFFR_X1 \registers_reg[3][5]  ( .D(n4016), .CK(n675), .RN(n6783), .Q(
        \registers[3][5] ), .QN(n4301) );
  DFFR_X1 \registers_reg[3][4]  ( .D(n4015), .CK(n675), .RN(n6786), .Q(
        \registers[3][4] ), .QN(n4300) );
  DFFR_X1 \registers_reg[3][3]  ( .D(n4014), .CK(n675), .RN(n6833), .Q(
        \registers[3][3] ), .QN(n4299) );
  DFFR_X1 \registers_reg[3][2]  ( .D(n4013), .CK(n675), .RN(n6775), .Q(
        \registers[3][2] ), .QN(n4298) );
  DFFR_X1 \registers_reg[3][1]  ( .D(n4012), .CK(n675), .RN(n6769), .Q(
        \registers[3][1] ), .QN(n4297) );
  DFFR_X1 \registers_reg[3][0]  ( .D(n4011), .CK(n675), .RN(n6856), .Q(
        \registers[3][0] ), .QN(n4296) );
  DFFR_X1 \registers_reg[4][31]  ( .D(n4010), .CK(n675), .RN(n6836), .Q(
        \registers[4][31] ) );
  DFFR_X1 \registers_reg[4][30]  ( .D(n4009), .CK(n675), .RN(n6830), .Q(
        \registers[4][30] ) );
  DFFR_X1 \registers_reg[4][29]  ( .D(n4008), .CK(n675), .RN(n6825), .Q(
        \registers[4][29] ) );
  DFFR_X1 \registers_reg[4][28]  ( .D(n4007), .CK(n675), .RN(n6819), .Q(
        \registers[4][28] ) );
  DFFR_X1 \registers_reg[4][27]  ( .D(n4006), .CK(n675), .RN(n6839), .Q(
        \registers[4][27] ) );
  DFFR_X1 \registers_reg[4][26]  ( .D(n4005), .CK(n675), .RN(n6811), .Q(
        \registers[4][26] ) );
  DFFR_X1 \registers_reg[4][25]  ( .D(n4004), .CK(n675), .RN(n6814), .Q(
        \registers[4][25] ) );
  DFFR_X1 \registers_reg[4][24]  ( .D(n4003), .CK(n675), .RN(n6806), .Q(
        \registers[4][24] ) );
  DFFR_X1 \registers_reg[4][23]  ( .D(n4002), .CK(n675), .RN(n6842), .Q(
        \registers[4][23] ) );
  DFFR_X1 \registers_reg[4][22]  ( .D(n4001), .CK(n675), .RN(n6794), .Q(
        \registers[4][22] ) );
  DFFR_X1 \registers_reg[4][21]  ( .D(n4000), .CK(n675), .RN(n6797), .Q(
        \registers[4][21] ) );
  DFFR_X1 \registers_reg[4][20]  ( .D(n3999), .CK(n675), .RN(n6789), .Q(
        \registers[4][20] ) );
  DFFR_X1 \registers_reg[4][19]  ( .D(n3998), .CK(n675), .RN(n6844), .Q(
        \registers[4][19] ) );
  DFFR_X1 \registers_reg[4][18]  ( .D(n3997), .CK(n675), .RN(n6778), .Q(
        \registers[4][18] ) );
  DFFR_X1 \registers_reg[4][17]  ( .D(n3996), .CK(n675), .RN(n6781), .Q(
        \registers[4][17] ) );
  DFFR_X1 \registers_reg[4][16]  ( .D(n3995), .CK(n675), .RN(n6772), .Q(
        \registers[4][16] ) );
  DFFR_X1 \registers_reg[4][15]  ( .D(n3994), .CK(n675), .RN(n6847), .Q(
        \registers[4][15] ) );
  DFFR_X1 \registers_reg[4][14]  ( .D(n3993), .CK(n675), .RN(n6828), .Q(
        \registers[4][14] ) );
  DFFR_X1 \registers_reg[4][13]  ( .D(n3992), .CK(n675), .RN(n6822), .Q(
        \registers[4][13] ) );
  DFFR_X1 \registers_reg[4][12]  ( .D(n3991), .CK(n675), .RN(n6817), .Q(
        \registers[4][12] ) );
  DFFR_X1 \registers_reg[4][11]  ( .D(n3990), .CK(n675), .RN(n6850), .Q(
        \registers[4][11] ) );
  DFFR_X1 \registers_reg[4][10]  ( .D(n3989), .CK(n675), .RN(n6808), .Q(
        \registers[4][10] ) );
  DFFR_X1 \registers_reg[4][9]  ( .D(n3988), .CK(n675), .RN(n6800), .Q(
        \registers[4][9] ) );
  DFFR_X1 \registers_reg[4][8]  ( .D(n3987), .CK(n675), .RN(n6803), .Q(
        \registers[4][8] ) );
  DFFR_X1 \registers_reg[4][7]  ( .D(n3986), .CK(n675), .RN(n6853), .Q(
        \registers[4][7] ) );
  DFFR_X1 \registers_reg[4][6]  ( .D(n3985), .CK(n675), .RN(n6792), .Q(
        \registers[4][6] ) );
  DFFR_X1 \registers_reg[4][5]  ( .D(n3984), .CK(n675), .RN(n6783), .Q(
        \registers[4][5] ) );
  DFFR_X1 \registers_reg[4][4]  ( .D(n3983), .CK(n675), .RN(n6786), .Q(
        \registers[4][4] ) );
  DFFR_X1 \registers_reg[4][3]  ( .D(n3982), .CK(n675), .RN(n6833), .Q(
        \registers[4][3] ) );
  DFFR_X1 \registers_reg[4][2]  ( .D(n3981), .CK(n675), .RN(n6775), .Q(
        \registers[4][2] ) );
  DFFR_X1 \registers_reg[4][1]  ( .D(n3980), .CK(n675), .RN(n6769), .Q(
        \registers[4][1] ) );
  DFFR_X1 \registers_reg[4][0]  ( .D(n3979), .CK(n675), .RN(n6856), .Q(
        \registers[4][0] ) );
  DFFR_X1 \registers_reg[5][31]  ( .D(n3978), .CK(n675), .RN(n6836), .Q(
        \registers[5][31] ) );
  DFFR_X1 \registers_reg[5][30]  ( .D(n3977), .CK(n675), .RN(n6830), .Q(
        \registers[5][30] ) );
  DFFR_X1 \registers_reg[5][29]  ( .D(n3976), .CK(n675), .RN(n6825), .Q(
        \registers[5][29] ) );
  DFFR_X1 \registers_reg[5][28]  ( .D(n3975), .CK(n675), .RN(n6819), .Q(
        \registers[5][28] ) );
  DFFR_X1 \registers_reg[5][27]  ( .D(n3974), .CK(n675), .RN(n6839), .Q(
        \registers[5][27] ) );
  DFFR_X1 \registers_reg[5][26]  ( .D(n3973), .CK(n675), .RN(n6811), .Q(
        \registers[5][26] ) );
  DFFR_X1 \registers_reg[5][25]  ( .D(n3972), .CK(n675), .RN(n6814), .Q(
        \registers[5][25] ) );
  DFFR_X1 \registers_reg[5][24]  ( .D(n3971), .CK(n675), .RN(n6805), .Q(
        \registers[5][24] ) );
  DFFR_X1 \registers_reg[5][23]  ( .D(n3970), .CK(n675), .RN(n6842), .Q(
        \registers[5][23] ) );
  DFFR_X1 \registers_reg[5][22]  ( .D(n3969), .CK(n675), .RN(n6794), .Q(
        \registers[5][22] ) );
  DFFR_X1 \registers_reg[5][21]  ( .D(n3968), .CK(n675), .RN(n6797), .Q(
        \registers[5][21] ) );
  DFFR_X1 \registers_reg[5][20]  ( .D(n3967), .CK(n675), .RN(n6789), .Q(
        \registers[5][20] ) );
  DFFR_X1 \registers_reg[5][19]  ( .D(n3966), .CK(n675), .RN(n6844), .Q(
        \registers[5][19] ) );
  DFFR_X1 \registers_reg[5][18]  ( .D(n3965), .CK(n675), .RN(n6778), .Q(
        \registers[5][18] ) );
  DFFR_X1 \registers_reg[5][17]  ( .D(n3964), .CK(n675), .RN(n6780), .Q(
        \registers[5][17] ) );
  DFFR_X1 \registers_reg[5][16]  ( .D(n3963), .CK(n675), .RN(n6772), .Q(
        \registers[5][16] ) );
  DFFR_X1 \registers_reg[5][15]  ( .D(n3962), .CK(n675), .RN(n6847), .Q(
        \registers[5][15] ) );
  DFFR_X1 \registers_reg[5][14]  ( .D(n3961), .CK(n675), .RN(n6828), .Q(
        \registers[5][14] ) );
  DFFR_X1 \registers_reg[5][13]  ( .D(n3960), .CK(n675), .RN(n6822), .Q(
        \registers[5][13] ) );
  DFFR_X1 \registers_reg[5][12]  ( .D(n3959), .CK(n675), .RN(n6817), .Q(
        \registers[5][12] ) );
  DFFR_X1 \registers_reg[5][11]  ( .D(n3958), .CK(n675), .RN(n6850), .Q(
        \registers[5][11] ) );
  DFFR_X1 \registers_reg[5][10]  ( .D(n3957), .CK(n675), .RN(n6808), .Q(
        \registers[5][10] ) );
  DFFR_X1 \registers_reg[5][9]  ( .D(n3956), .CK(n675), .RN(n6800), .Q(
        \registers[5][9] ) );
  DFFR_X1 \registers_reg[5][8]  ( .D(n3955), .CK(n675), .RN(n6803), .Q(
        \registers[5][8] ) );
  DFFR_X1 \registers_reg[5][7]  ( .D(n3954), .CK(n675), .RN(n6853), .Q(
        \registers[5][7] ) );
  DFFR_X1 \registers_reg[5][6]  ( .D(n3953), .CK(n675), .RN(n6792), .Q(
        \registers[5][6] ) );
  DFFR_X1 \registers_reg[5][5]  ( .D(n3952), .CK(n675), .RN(n6783), .Q(
        \registers[5][5] ) );
  DFFR_X1 \registers_reg[5][4]  ( .D(n3951), .CK(n675), .RN(n6786), .Q(
        \registers[5][4] ) );
  DFFR_X1 \registers_reg[5][3]  ( .D(n3950), .CK(n675), .RN(n6833), .Q(
        \registers[5][3] ) );
  DFFR_X1 \registers_reg[5][2]  ( .D(n3949), .CK(n675), .RN(n6775), .Q(
        \registers[5][2] ) );
  DFFR_X1 \registers_reg[5][1]  ( .D(n3948), .CK(n675), .RN(n6769), .Q(
        \registers[5][1] ) );
  DFFR_X1 \registers_reg[5][0]  ( .D(n3947), .CK(n675), .RN(n6856), .Q(
        \registers[5][0] ) );
  DFFR_X1 \registers_reg[6][31]  ( .D(n3946), .CK(n675), .RN(n6836), .Q(
        \registers[6][31] ) );
  DFFR_X1 \registers_reg[6][30]  ( .D(n3945), .CK(n675), .RN(n6830), .Q(
        \registers[6][30] ) );
  DFFR_X1 \registers_reg[6][29]  ( .D(n3944), .CK(n675), .RN(n6825), .Q(
        \registers[6][29] ) );
  DFFR_X1 \registers_reg[6][28]  ( .D(n3943), .CK(n675), .RN(n6819), .Q(
        \registers[6][28] ) );
  DFFR_X1 \registers_reg[6][27]  ( .D(n3942), .CK(n675), .RN(n6839), .Q(
        \registers[6][27] ) );
  DFFR_X1 \registers_reg[6][26]  ( .D(n3941), .CK(n675), .RN(n6811), .Q(
        \registers[6][26] ) );
  DFFR_X1 \registers_reg[6][25]  ( .D(n3940), .CK(n675), .RN(n6814), .Q(
        \registers[6][25] ) );
  DFFR_X1 \registers_reg[6][24]  ( .D(n3939), .CK(n675), .RN(n6805), .Q(
        \registers[6][24] ) );
  DFFR_X1 \registers_reg[6][23]  ( .D(n3938), .CK(n675), .RN(n6841), .Q(
        \registers[6][23] ) );
  DFFR_X1 \registers_reg[6][22]  ( .D(n3937), .CK(n675), .RN(n6794), .Q(
        \registers[6][22] ) );
  DFFR_X1 \registers_reg[6][21]  ( .D(n3936), .CK(n675), .RN(n6797), .Q(
        \registers[6][21] ) );
  DFFR_X1 \registers_reg[6][20]  ( .D(n3935), .CK(n675), .RN(n6789), .Q(
        \registers[6][20] ) );
  DFFR_X1 \registers_reg[6][19]  ( .D(n3934), .CK(n675), .RN(n6844), .Q(
        \registers[6][19] ) );
  DFFR_X1 \registers_reg[6][18]  ( .D(n3933), .CK(n675), .RN(n6778), .Q(
        \registers[6][18] ) );
  DFFR_X1 \registers_reg[6][17]  ( .D(n3932), .CK(n675), .RN(n6780), .Q(
        \registers[6][17] ) );
  DFFR_X1 \registers_reg[6][16]  ( .D(n3931), .CK(n675), .RN(n6772), .Q(
        \registers[6][16] ) );
  DFFR_X1 \registers_reg[6][15]  ( .D(n3930), .CK(n675), .RN(n6847), .Q(
        \registers[6][15] ) );
  DFFR_X1 \registers_reg[6][14]  ( .D(n3929), .CK(n675), .RN(n6827), .Q(
        \registers[6][14] ) );
  DFFR_X1 \registers_reg[6][13]  ( .D(n3928), .CK(n675), .RN(n6822), .Q(
        \registers[6][13] ) );
  DFFR_X1 \registers_reg[6][12]  ( .D(n3927), .CK(n675), .RN(n6816), .Q(
        \registers[6][12] ) );
  DFFR_X1 \registers_reg[6][11]  ( .D(n3926), .CK(n675), .RN(n6850), .Q(
        \registers[6][11] ) );
  DFFR_X1 \registers_reg[6][10]  ( .D(n3925), .CK(n675), .RN(n6808), .Q(
        \registers[6][10] ) );
  DFFR_X1 \registers_reg[6][9]  ( .D(n3924), .CK(n675), .RN(n6800), .Q(
        \registers[6][9] ) );
  DFFR_X1 \registers_reg[6][8]  ( .D(n3923), .CK(n675), .RN(n6803), .Q(
        \registers[6][8] ) );
  DFFR_X1 \registers_reg[6][7]  ( .D(n3922), .CK(n675), .RN(n6853), .Q(
        \registers[6][7] ) );
  DFFR_X1 \registers_reg[6][6]  ( .D(n3921), .CK(n675), .RN(n6791), .Q(
        \registers[6][6] ) );
  DFFR_X1 \registers_reg[6][5]  ( .D(n3920), .CK(n675), .RN(n6783), .Q(
        \registers[6][5] ) );
  DFFR_X1 \registers_reg[6][4]  ( .D(n3919), .CK(n675), .RN(n6786), .Q(
        \registers[6][4] ) );
  DFFR_X1 \registers_reg[6][3]  ( .D(n3918), .CK(n675), .RN(n6833), .Q(
        \registers[6][3] ) );
  DFFR_X1 \registers_reg[6][2]  ( .D(n3917), .CK(n675), .RN(n6775), .Q(
        \registers[6][2] ) );
  DFFR_X1 \registers_reg[6][1]  ( .D(n3916), .CK(n675), .RN(n6769), .Q(
        \registers[6][1] ) );
  DFFR_X1 \registers_reg[6][0]  ( .D(n3915), .CK(n675), .RN(n6856), .Q(
        \registers[6][0] ) );
  DFFR_X1 \registers_reg[7][31]  ( .D(n3914), .CK(n675), .RN(n6836), .Q(
        \registers[7][31] ) );
  DFFR_X1 \registers_reg[7][30]  ( .D(n3913), .CK(n675), .RN(n6830), .Q(
        \registers[7][30] ) );
  DFFR_X1 \registers_reg[7][29]  ( .D(n3912), .CK(n675), .RN(n6825), .Q(
        \registers[7][29] ) );
  DFFR_X1 \registers_reg[7][28]  ( .D(n3911), .CK(n675), .RN(n6819), .Q(
        \registers[7][28] ) );
  DFFR_X1 \registers_reg[7][27]  ( .D(n3910), .CK(n675), .RN(n6839), .Q(
        \registers[7][27] ) );
  DFFR_X1 \registers_reg[7][26]  ( .D(n3909), .CK(n675), .RN(n6811), .Q(
        \registers[7][26] ) );
  DFFR_X1 \registers_reg[7][25]  ( .D(n3908), .CK(n675), .RN(n6814), .Q(
        \registers[7][25] ) );
  DFFR_X1 \registers_reg[7][24]  ( .D(n3907), .CK(n675), .RN(n6805), .Q(
        \registers[7][24] ) );
  DFFR_X1 \registers_reg[7][23]  ( .D(n3906), .CK(n675), .RN(n6841), .Q(
        \registers[7][23] ) );
  DFFR_X1 \registers_reg[7][22]  ( .D(n3905), .CK(n675), .RN(n6794), .Q(
        \registers[7][22] ) );
  DFFR_X1 \registers_reg[7][21]  ( .D(n3904), .CK(n675), .RN(n6797), .Q(
        \registers[7][21] ) );
  DFFR_X1 \registers_reg[7][20]  ( .D(n3903), .CK(n675), .RN(n6789), .Q(
        \registers[7][20] ) );
  DFFR_X1 \registers_reg[7][19]  ( .D(n3902), .CK(n675), .RN(n6844), .Q(
        \registers[7][19] ) );
  DFFR_X1 \registers_reg[7][18]  ( .D(n3901), .CK(n675), .RN(n6777), .Q(
        \registers[7][18] ) );
  DFFR_X1 \registers_reg[7][17]  ( .D(n3900), .CK(n675), .RN(n6780), .Q(
        \registers[7][17] ) );
  DFFR_X1 \registers_reg[7][16]  ( .D(n3899), .CK(n675), .RN(n6772), .Q(
        \registers[7][16] ) );
  DFFR_X1 \registers_reg[7][15]  ( .D(n3898), .CK(n675), .RN(n6847), .Q(
        \registers[7][15] ) );
  DFFR_X1 \registers_reg[7][14]  ( .D(n3897), .CK(n675), .RN(n6827), .Q(
        \registers[7][14] ) );
  DFFR_X1 \registers_reg[7][13]  ( .D(n3896), .CK(n675), .RN(n6822), .Q(
        \registers[7][13] ) );
  DFFR_X1 \registers_reg[7][12]  ( .D(n3895), .CK(n675), .RN(n6816), .Q(
        \registers[7][12] ) );
  DFFR_X1 \registers_reg[7][11]  ( .D(n3894), .CK(n675), .RN(n6850), .Q(
        \registers[7][11] ) );
  DFFR_X1 \registers_reg[7][10]  ( .D(n3893), .CK(n675), .RN(n6808), .Q(
        \registers[7][10] ) );
  DFFR_X1 \registers_reg[7][9]  ( .D(n3892), .CK(n675), .RN(n6800), .Q(
        \registers[7][9] ) );
  DFFR_X1 \registers_reg[7][8]  ( .D(n3891), .CK(n675), .RN(n6803), .Q(
        \registers[7][8] ) );
  DFFR_X1 \registers_reg[7][7]  ( .D(n3890), .CK(n675), .RN(n6853), .Q(
        \registers[7][7] ) );
  DFFR_X1 \registers_reg[7][6]  ( .D(n3889), .CK(n675), .RN(n6791), .Q(
        \registers[7][6] ) );
  DFFR_X1 \registers_reg[7][5]  ( .D(n3888), .CK(n675), .RN(n6783), .Q(
        \registers[7][5] ) );
  DFFR_X1 \registers_reg[7][4]  ( .D(n3887), .CK(n675), .RN(n6786), .Q(
        \registers[7][4] ) );
  DFFR_X1 \registers_reg[7][3]  ( .D(n3886), .CK(n675), .RN(n6833), .Q(
        \registers[7][3] ) );
  DFFR_X1 \registers_reg[7][2]  ( .D(n3885), .CK(n675), .RN(n6775), .Q(
        \registers[7][2] ) );
  DFFR_X1 \registers_reg[7][1]  ( .D(n3884), .CK(n675), .RN(n6769), .Q(
        \registers[7][1] ) );
  DFFR_X1 \registers_reg[7][0]  ( .D(n3883), .CK(n675), .RN(n6856), .Q(
        \registers[7][0] ) );
  DFFR_X1 \registers_reg[8][31]  ( .D(n3882), .CK(n675), .RN(n6836), .Q(
        \registers[8][31] ), .QN(n5840) );
  DFFR_X1 \registers_reg[8][30]  ( .D(n3881), .CK(n675), .RN(n6830), .Q(
        \registers[8][30] ), .QN(n5838) );
  DFFR_X1 \registers_reg[8][29]  ( .D(n3880), .CK(n675), .RN(n6825), .Q(
        \registers[8][29] ), .QN(n5836) );
  DFFR_X1 \registers_reg[8][28]  ( .D(n3879), .CK(n675), .RN(n6819), .Q(
        \registers[8][28] ), .QN(n5834) );
  DFFR_X1 \registers_reg[8][27]  ( .D(n3878), .CK(n675), .RN(n6838), .Q(
        \registers[8][27] ), .QN(n5833) );
  DFFR_X1 \registers_reg[8][26]  ( .D(n3877), .CK(n675), .RN(n6811), .Q(
        \registers[8][26] ), .QN(n5832) );
  DFFR_X1 \registers_reg[8][25]  ( .D(n3876), .CK(n675), .RN(n6814), .Q(
        \registers[8][25] ), .QN(n5831) );
  DFFR_X1 \registers_reg[8][24]  ( .D(n3875), .CK(n675), .RN(n6805), .Q(
        \registers[8][24] ), .QN(n5830) );
  DFFR_X1 \registers_reg[8][23]  ( .D(n3874), .CK(n675), .RN(n6841), .Q(
        \registers[8][23] ), .QN(n5829) );
  DFFR_X1 \registers_reg[8][22]  ( .D(n3873), .CK(n675), .RN(n6794), .Q(
        \registers[8][22] ), .QN(n5828) );
  DFFR_X1 \registers_reg[8][21]  ( .D(n3872), .CK(n675), .RN(n6797), .Q(
        \registers[8][21] ), .QN(n5826) );
  DFFR_X1 \registers_reg[8][20]  ( .D(n3871), .CK(n675), .RN(n6789), .Q(
        \registers[8][20] ), .QN(n5824) );
  DFFR_X1 \registers_reg[8][19]  ( .D(n3870), .CK(n675), .RN(n6844), .Q(
        \registers[8][19] ), .QN(n5822) );
  DFFR_X1 \registers_reg[8][18]  ( .D(n3869), .CK(n675), .RN(n6777), .Q(
        \registers[8][18] ), .QN(n5820) );
  DFFR_X1 \registers_reg[8][17]  ( .D(n3868), .CK(n675), .RN(n6780), .Q(
        \registers[8][17] ), .QN(n5818) );
  DFFR_X1 \registers_reg[8][16]  ( .D(n3867), .CK(n675), .RN(n6772), .Q(
        \registers[8][16] ), .QN(n5816) );
  DFFR_X1 \registers_reg[8][15]  ( .D(n3866), .CK(n675), .RN(n6847), .Q(
        \registers[8][15] ), .QN(n5814) );
  DFFR_X1 \registers_reg[8][14]  ( .D(n3865), .CK(n675), .RN(n6827), .Q(
        \registers[8][14] ), .QN(n5812) );
  DFFR_X1 \registers_reg[8][13]  ( .D(n3864), .CK(n675), .RN(n6822), .Q(
        \registers[8][13] ), .QN(n5810) );
  DFFR_X1 \registers_reg[8][12]  ( .D(n3863), .CK(n675), .RN(n6816), .Q(
        \registers[8][12] ), .QN(n5808) );
  DFFR_X1 \registers_reg[8][11]  ( .D(n3862), .CK(n675), .RN(n6850), .Q(
        \registers[8][11] ), .QN(n5806) );
  DFFR_X1 \registers_reg[8][10]  ( .D(n3861), .CK(n675), .RN(n6808), .Q(
        \registers[8][10] ), .QN(n5804) );
  DFFR_X1 \registers_reg[8][9]  ( .D(n3860), .CK(n675), .RN(n6800), .Q(
        \registers[8][9] ), .QN(n5802) );
  DFFR_X1 \registers_reg[8][8]  ( .D(n3859), .CK(n675), .RN(n6802), .Q(
        \registers[8][8] ), .QN(n5800) );
  DFFR_X1 \registers_reg[8][7]  ( .D(n3858), .CK(n675), .RN(n6853), .Q(
        \registers[8][7] ), .QN(n5798) );
  DFFR_X1 \registers_reg[8][6]  ( .D(n3857), .CK(n675), .RN(n6791), .Q(
        \registers[8][6] ), .QN(n5796) );
  DFFR_X1 \registers_reg[8][5]  ( .D(n3856), .CK(n675), .RN(n6783), .Q(
        \registers[8][5] ), .QN(n5794) );
  DFFR_X1 \registers_reg[8][4]  ( .D(n3855), .CK(n675), .RN(n6786), .Q(
        \registers[8][4] ), .QN(n5792) );
  DFFR_X1 \registers_reg[8][3]  ( .D(n3854), .CK(n675), .RN(n6833), .Q(
        \registers[8][3] ), .QN(n5790) );
  DFFR_X1 \registers_reg[8][2]  ( .D(n3853), .CK(n675), .RN(n6775), .Q(
        \registers[8][2] ), .QN(n5788) );
  DFFR_X1 \registers_reg[8][1]  ( .D(n3852), .CK(n675), .RN(n6769), .Q(
        \registers[8][1] ), .QN(n5786) );
  DFFR_X1 \registers_reg[8][0]  ( .D(n3851), .CK(n675), .RN(n6855), .Q(
        \registers[8][0] ), .QN(n5784) );
  DFFR_X1 \registers_reg[9][31]  ( .D(n3850), .CK(n675), .RN(n6836), .Q(
        \registers[9][31] ), .QN(n2850) );
  DFFR_X1 \registers_reg[9][30]  ( .D(n3849), .CK(n675), .RN(n6830), .Q(
        \registers[9][30] ), .QN(n2848) );
  DFFR_X1 \registers_reg[9][29]  ( .D(n3848), .CK(n675), .RN(n6824), .Q(
        \registers[9][29] ), .QN(n2846) );
  DFFR_X1 \registers_reg[9][28]  ( .D(n3847), .CK(n675), .RN(n6819), .Q(
        \registers[9][28] ), .QN(n2844) );
  DFFR_X1 \registers_reg[9][27]  ( .D(n3846), .CK(n675), .RN(n6838), .Q(
        \registers[9][27] ), .QN(n2843) );
  DFFR_X1 \registers_reg[9][26]  ( .D(n3845), .CK(n675), .RN(n6811), .Q(
        \registers[9][26] ), .QN(n2842) );
  DFFR_X1 \registers_reg[9][25]  ( .D(n3844), .CK(n675), .RN(n6813), .Q(
        \registers[9][25] ), .QN(n2841) );
  DFFR_X1 \registers_reg[9][24]  ( .D(n3843), .CK(n675), .RN(n6805), .Q(
        \registers[9][24] ), .QN(n2840) );
  DFFR_X1 \registers_reg[9][23]  ( .D(n3842), .CK(n675), .RN(n6841), .Q(
        \registers[9][23] ), .QN(n2839) );
  DFFR_X1 \registers_reg[9][22]  ( .D(n3841), .CK(n675), .RN(n6794), .Q(
        \registers[9][22] ), .QN(n2838) );
  DFFR_X1 \registers_reg[9][21]  ( .D(n3840), .CK(n675), .RN(n6797), .Q(
        \registers[9][21] ), .QN(n2836) );
  DFFR_X1 \registers_reg[9][20]  ( .D(n3839), .CK(n675), .RN(n6788), .Q(
        \registers[9][20] ), .QN(n2834) );
  DFFR_X1 \registers_reg[9][19]  ( .D(n3838), .CK(n675), .RN(n6844), .Q(
        \registers[9][19] ), .QN(n2832) );
  DFFR_X1 \registers_reg[9][18]  ( .D(n3837), .CK(n675), .RN(n6777), .Q(
        \registers[9][18] ), .QN(n2830) );
  DFFR_X1 \registers_reg[9][17]  ( .D(n3836), .CK(n675), .RN(n6780), .Q(
        \registers[9][17] ), .QN(n2828) );
  DFFR_X1 \registers_reg[9][16]  ( .D(n3835), .CK(n675), .RN(n6772), .Q(
        \registers[9][16] ), .QN(n2826) );
  DFFR_X1 \registers_reg[9][15]  ( .D(n3834), .CK(n675), .RN(n6847), .Q(
        \registers[9][15] ), .QN(n2822) );
  DFFR_X1 \registers_reg[9][14]  ( .D(n3833), .CK(n675), .RN(n6827), .Q(
        \registers[9][14] ), .QN(n2820) );
  DFFR_X1 \registers_reg[9][13]  ( .D(n3832), .CK(n675), .RN(n6822), .Q(
        \registers[9][13] ), .QN(n2818) );
  DFFR_X1 \registers_reg[9][12]  ( .D(n3831), .CK(n675), .RN(n6816), .Q(
        \registers[9][12] ), .QN(n2816) );
  DFFR_X1 \registers_reg[9][11]  ( .D(n3830), .CK(n675), .RN(n6850), .Q(
        \registers[9][11] ), .QN(n2814) );
  DFFR_X1 \registers_reg[9][10]  ( .D(n3829), .CK(n675), .RN(n6808), .Q(
        \registers[9][10] ), .QN(n2812) );
  DFFR_X1 \registers_reg[9][9]  ( .D(n3828), .CK(n675), .RN(n6800), .Q(
        \registers[9][9] ), .QN(n2810) );
  DFFR_X1 \registers_reg[9][8]  ( .D(n3827), .CK(n675), .RN(n6802), .Q(
        \registers[9][8] ), .QN(n2808) );
  DFFR_X1 \registers_reg[9][7]  ( .D(n3826), .CK(n675), .RN(n6853), .Q(
        \registers[9][7] ), .QN(n2806) );
  DFFR_X1 \registers_reg[9][6]  ( .D(n3825), .CK(n675), .RN(n6791), .Q(
        \registers[9][6] ), .QN(n2804) );
  DFFR_X1 \registers_reg[9][5]  ( .D(n3824), .CK(n675), .RN(n6783), .Q(
        \registers[9][5] ), .QN(n2802) );
  DFFR_X1 \registers_reg[9][4]  ( .D(n3823), .CK(n675), .RN(n6786), .Q(
        \registers[9][4] ), .QN(n2800) );
  DFFR_X1 \registers_reg[9][3]  ( .D(n3822), .CK(n675), .RN(n6833), .Q(
        \registers[9][3] ), .QN(n2798) );
  DFFR_X1 \registers_reg[9][2]  ( .D(n3821), .CK(n675), .RN(n6775), .Q(
        \registers[9][2] ), .QN(n2796) );
  DFFR_X1 \registers_reg[9][1]  ( .D(n3820), .CK(n675), .RN(n6769), .Q(
        \registers[9][1] ), .QN(n2794) );
  DFFR_X1 \registers_reg[9][0]  ( .D(n3819), .CK(n675), .RN(n6855), .Q(
        \registers[9][0] ), .QN(n2792) );
  DFFR_X1 \registers_reg[10][31]  ( .D(n3818), .CK(n675), .RN(n6835), .Q(
        \registers[10][31] ), .QN(n4346) );
  DFFR_X1 \registers_reg[10][30]  ( .D(n3817), .CK(n675), .RN(n6830), .Q(
        \registers[10][30] ), .QN(n4345) );
  DFFR_X1 \registers_reg[10][29]  ( .D(n3816), .CK(n675), .RN(n6824), .Q(
        \registers[10][29] ), .QN(n5773) );
  DFFR_X1 \registers_reg[10][28]  ( .D(n3815), .CK(n675), .RN(n6819), .Q(
        \registers[10][28] ), .QN(n4344) );
  DFFR_X1 \registers_reg[10][27]  ( .D(n3814), .CK(n675), .RN(n6838), .Q(
        \registers[10][27] ), .QN(n4343) );
  DFFR_X1 \registers_reg[10][26]  ( .D(n3813), .CK(n675), .RN(n6811), .Q(
        \registers[10][26] ), .QN(n5772) );
  DFFR_X1 \registers_reg[10][25]  ( .D(n3812), .CK(n675), .RN(n6813), .Q(
        \registers[10][25] ), .QN(n4342) );
  DFFR_X1 \registers_reg[10][24]  ( .D(n3811), .CK(n675), .RN(n6805), .Q(
        \registers[10][24] ), .QN(n4341) );
  DFFR_X1 \registers_reg[10][23]  ( .D(n3810), .CK(n675), .RN(n6841), .Q(
        \registers[10][23] ), .QN(n5771) );
  DFFR_X1 \registers_reg[10][22]  ( .D(n3809), .CK(n675), .RN(n6794), .Q(
        \registers[10][22] ), .QN(n4340) );
  DFFR_X1 \registers_reg[10][21]  ( .D(n3808), .CK(n675), .RN(n6797), .Q(
        \registers[10][21] ), .QN(n4339) );
  DFFR_X1 \registers_reg[10][20]  ( .D(n3807), .CK(n675), .RN(n6788), .Q(
        \registers[10][20] ), .QN(n5770) );
  DFFR_X1 \registers_reg[10][19]  ( .D(n3806), .CK(n675), .RN(n6844), .Q(
        \registers[10][19] ), .QN(n4338) );
  DFFR_X1 \registers_reg[10][18]  ( .D(n3805), .CK(n675), .RN(n6777), .Q(
        \registers[10][18] ), .QN(n4337) );
  DFFR_X1 \registers_reg[10][17]  ( .D(n3804), .CK(n675), .RN(n6780), .Q(
        \registers[10][17] ), .QN(n5769) );
  DFFR_X1 \registers_reg[10][16]  ( .D(n3803), .CK(n675), .RN(n6772), .Q(
        \registers[10][16] ), .QN(n4336) );
  DFFR_X1 \registers_reg[10][15]  ( .D(n3802), .CK(n675), .RN(n6847), .Q(
        \registers[10][15] ), .QN(n4335) );
  DFFR_X1 \registers_reg[10][14]  ( .D(n3801), .CK(n675), .RN(n6827), .Q(
        \registers[10][14] ), .QN(n5768) );
  DFFR_X1 \registers_reg[10][13]  ( .D(n3800), .CK(n675), .RN(n6822), .Q(
        \registers[10][13] ), .QN(n4334) );
  DFFR_X1 \registers_reg[10][12]  ( .D(n3799), .CK(n675), .RN(n6816), .Q(
        \registers[10][12] ), .QN(n4333) );
  DFFR_X1 \registers_reg[10][11]  ( .D(n3798), .CK(n675), .RN(n6850), .Q(
        \registers[10][11] ), .QN(n5767) );
  DFFR_X1 \registers_reg[10][10]  ( .D(n3797), .CK(n675), .RN(n6808), .Q(
        \registers[10][10] ), .QN(n4332) );
  DFFR_X1 \registers_reg[10][9]  ( .D(n3796), .CK(n675), .RN(n6799), .Q(
        \registers[10][9] ), .QN(n4331) );
  DFFR_X1 \registers_reg[10][8]  ( .D(n3795), .CK(n675), .RN(n6802), .Q(
        \registers[10][8] ), .QN(n5766) );
  DFFR_X1 \registers_reg[10][7]  ( .D(n3794), .CK(n675), .RN(n6852), .Q(
        \registers[10][7] ), .QN(n4330) );
  DFFR_X1 \registers_reg[10][6]  ( .D(n3793), .CK(n675), .RN(n6791), .Q(
        \registers[10][6] ), .QN(n4329) );
  DFFR_X1 \registers_reg[10][5]  ( .D(n3792), .CK(n675), .RN(n6783), .Q(
        \registers[10][5] ), .QN(n5765) );
  DFFR_X1 \registers_reg[10][4]  ( .D(n3791), .CK(n675), .RN(n6786), .Q(
        \registers[10][4] ), .QN(n4328) );
  DFFR_X1 \registers_reg[10][3]  ( .D(n3790), .CK(n675), .RN(n6833), .Q(
        \registers[10][3] ), .QN(n4327) );
  DFFR_X1 \registers_reg[10][2]  ( .D(n3789), .CK(n675), .RN(n6774), .Q(
        \registers[10][2] ), .QN(n5764) );
  DFFR_X1 \registers_reg[10][1]  ( .D(n3788), .CK(n675), .RN(n6769), .Q(
        \registers[10][1] ), .QN(n4326) );
  DFFR_X1 \registers_reg[10][0]  ( .D(n3787), .CK(n675), .RN(n6855), .Q(
        \registers[10][0] ), .QN(n4325) );
  DFFR_X1 \registers_reg[11][31]  ( .D(n3786), .CK(n675), .RN(n6835), .Q(
        \registers[11][31] ), .QN(n2753) );
  DFFR_X1 \registers_reg[11][30]  ( .D(n3785), .CK(n675), .RN(n6830), .Q(
        \registers[11][30] ), .QN(n2752) );
  DFFR_X1 \registers_reg[11][29]  ( .D(n3784), .CK(n675), .RN(n6824), .Q(
        \registers[11][29] ), .QN(n2780) );
  DFFR_X1 \registers_reg[11][28]  ( .D(n3783), .CK(n675), .RN(n6819), .Q(
        \registers[11][28] ), .QN(n2751) );
  DFFR_X1 \registers_reg[11][27]  ( .D(n3782), .CK(n675), .RN(n6838), .Q(
        \registers[11][27] ), .QN(n2750) );
  DFFR_X1 \registers_reg[11][26]  ( .D(n3781), .CK(n675), .RN(n6810), .Q(
        \registers[11][26] ), .QN(n2779) );
  DFFR_X1 \registers_reg[11][25]  ( .D(n3780), .CK(n675), .RN(n6813), .Q(
        \registers[11][25] ), .QN(n2749) );
  DFFR_X1 \registers_reg[11][24]  ( .D(n3779), .CK(n675), .RN(n6805), .Q(
        \registers[11][24] ), .QN(n2748) );
  DFFR_X1 \registers_reg[11][23]  ( .D(n3778), .CK(n675), .RN(n6841), .Q(
        \registers[11][23] ), .QN(n2778) );
  DFFR_X1 \registers_reg[11][22]  ( .D(n3777), .CK(n675), .RN(n6794), .Q(
        \registers[11][22] ), .QN(n2747) );
  DFFR_X1 \registers_reg[11][21]  ( .D(n3776), .CK(n675), .RN(n6797), .Q(
        \registers[11][21] ), .QN(n2746) );
  DFFR_X1 \registers_reg[11][20]  ( .D(n3775), .CK(n675), .RN(n6788), .Q(
        \registers[11][20] ), .QN(n2777) );
  DFFR_X1 \registers_reg[11][19]  ( .D(n3774), .CK(n675), .RN(n6844), .Q(
        \registers[11][19] ), .QN(n2745) );
  DFFR_X1 \registers_reg[11][18]  ( .D(n3773), .CK(n675), .RN(n6777), .Q(
        \registers[11][18] ), .QN(n2744) );
  DFFR_X1 \registers_reg[11][17]  ( .D(n3772), .CK(n675), .RN(n6780), .Q(
        \registers[11][17] ), .QN(n2776) );
  DFFR_X1 \registers_reg[11][16]  ( .D(n3771), .CK(n675), .RN(n6772), .Q(
        \registers[11][16] ), .QN(n2743) );
  DFFR_X1 \registers_reg[11][15]  ( .D(n3770), .CK(n675), .RN(n6847), .Q(
        \registers[11][15] ), .QN(n2742) );
  DFFR_X1 \registers_reg[11][14]  ( .D(n3769), .CK(n675), .RN(n6827), .Q(
        \registers[11][14] ), .QN(n2775) );
  DFFR_X1 \registers_reg[11][13]  ( .D(n3768), .CK(n675), .RN(n6822), .Q(
        \registers[11][13] ), .QN(n2741) );
  DFFR_X1 \registers_reg[11][12]  ( .D(n3767), .CK(n675), .RN(n6816), .Q(
        \registers[11][12] ), .QN(n2740) );
  DFFR_X1 \registers_reg[11][11]  ( .D(n3766), .CK(n675), .RN(n6850), .Q(
        \registers[11][11] ), .QN(n2774) );
  DFFR_X1 \registers_reg[11][10]  ( .D(n3765), .CK(n675), .RN(n6808), .Q(
        \registers[11][10] ), .QN(n2739) );
  DFFR_X1 \registers_reg[11][9]  ( .D(n3764), .CK(n675), .RN(n6799), .Q(
        \registers[11][9] ), .QN(n2738) );
  DFFR_X1 \registers_reg[11][8]  ( .D(n3763), .CK(n675), .RN(n6802), .Q(
        \registers[11][8] ), .QN(n2773) );
  DFFR_X1 \registers_reg[11][7]  ( .D(n3762), .CK(n675), .RN(n6852), .Q(
        \registers[11][7] ), .QN(n2737) );
  DFFR_X1 \registers_reg[11][6]  ( .D(n3761), .CK(n675), .RN(n6791), .Q(
        \registers[11][6] ), .QN(n2736) );
  DFFR_X1 \registers_reg[11][5]  ( .D(n3760), .CK(n675), .RN(n6783), .Q(
        \registers[11][5] ), .QN(n2772) );
  DFFR_X1 \registers_reg[11][4]  ( .D(n3759), .CK(n675), .RN(n6786), .Q(
        \registers[11][4] ), .QN(n2735) );
  DFFR_X1 \registers_reg[11][3]  ( .D(n3758), .CK(n675), .RN(n6833), .Q(
        \registers[11][3] ), .QN(n2734) );
  DFFR_X1 \registers_reg[11][2]  ( .D(n3757), .CK(n675), .RN(n6774), .Q(
        \registers[11][2] ), .QN(n2771) );
  DFFR_X1 \registers_reg[11][1]  ( .D(n3756), .CK(n675), .RN(n6769), .Q(
        \registers[11][1] ), .QN(n2733) );
  DFFR_X1 \registers_reg[11][0]  ( .D(n3755), .CK(n675), .RN(n6855), .Q(
        \registers[11][0] ), .QN(n2732) );
  DFFR_X1 \registers_reg[12][31]  ( .D(n3754), .CK(n675), .RN(n6835), .Q(
        \registers[12][31] ) );
  DFFR_X1 \registers_reg[12][30]  ( .D(n3753), .CK(n675), .RN(n6830), .Q(
        \registers[12][30] ) );
  DFFR_X1 \registers_reg[12][29]  ( .D(n3752), .CK(n675), .RN(n6824), .Q(
        \registers[12][29] ) );
  DFFR_X1 \registers_reg[12][28]  ( .D(n3751), .CK(n675), .RN(n6819), .Q(
        \registers[12][28] ) );
  DFFR_X1 \registers_reg[12][27]  ( .D(n3750), .CK(n675), .RN(n6838), .Q(
        \registers[12][27] ) );
  DFFR_X1 \registers_reg[12][26]  ( .D(n3749), .CK(n675), .RN(n6810), .Q(
        \registers[12][26] ) );
  DFFR_X1 \registers_reg[12][25]  ( .D(n3748), .CK(n675), .RN(n6813), .Q(
        \registers[12][25] ) );
  DFFR_X1 \registers_reg[12][24]  ( .D(n3747), .CK(n675), .RN(n6805), .Q(
        \registers[12][24] ) );
  DFFR_X1 \registers_reg[12][23]  ( .D(n3746), .CK(n675), .RN(n6841), .Q(
        \registers[12][23] ) );
  DFFR_X1 \registers_reg[12][22]  ( .D(n3745), .CK(n675), .RN(n6794), .Q(
        \registers[12][22] ) );
  DFFR_X1 \registers_reg[12][21]  ( .D(n3744), .CK(n675), .RN(n6797), .Q(
        \registers[12][21] ) );
  DFFR_X1 \registers_reg[12][20]  ( .D(n3743), .CK(n675), .RN(n6788), .Q(
        \registers[12][20] ) );
  DFFR_X1 \registers_reg[12][19]  ( .D(n3742), .CK(n675), .RN(n6844), .Q(
        \registers[12][19] ) );
  DFFR_X1 \registers_reg[12][18]  ( .D(n3741), .CK(n675), .RN(n6777), .Q(
        \registers[12][18] ) );
  DFFR_X1 \registers_reg[12][17]  ( .D(n3740), .CK(n675), .RN(n6780), .Q(
        \registers[12][17] ) );
  DFFR_X1 \registers_reg[12][16]  ( .D(n3739), .CK(n675), .RN(n6771), .Q(
        \registers[12][16] ) );
  DFFR_X1 \registers_reg[12][15]  ( .D(n3738), .CK(n675), .RN(n6847), .Q(
        \registers[12][15] ) );
  DFFR_X1 \registers_reg[12][14]  ( .D(n3737), .CK(n675), .RN(n6827), .Q(
        \registers[12][14] ) );
  DFFR_X1 \registers_reg[12][13]  ( .D(n3736), .CK(n675), .RN(n6821), .Q(
        \registers[12][13] ) );
  DFFR_X1 \registers_reg[12][12]  ( .D(n3735), .CK(n675), .RN(n6816), .Q(
        \registers[12][12] ) );
  DFFR_X1 \registers_reg[12][11]  ( .D(n3734), .CK(n675), .RN(n6849), .Q(
        \registers[12][11] ) );
  DFFR_X1 \registers_reg[12][10]  ( .D(n3733), .CK(n675), .RN(n6808), .Q(
        \registers[12][10] ) );
  DFFR_X1 \registers_reg[12][9]  ( .D(n3732), .CK(n675), .RN(n6799), .Q(
        \registers[12][9] ) );
  DFFR_X1 \registers_reg[12][8]  ( .D(n3731), .CK(n675), .RN(n6802), .Q(
        \registers[12][8] ) );
  DFFR_X1 \registers_reg[12][7]  ( .D(n3730), .CK(n675), .RN(n6852), .Q(
        \registers[12][7] ) );
  DFFR_X1 \registers_reg[12][6]  ( .D(n3729), .CK(n675), .RN(n6791), .Q(
        \registers[12][6] ) );
  DFFR_X1 \registers_reg[12][5]  ( .D(n3728), .CK(n675), .RN(n6783), .Q(
        \registers[12][5] ) );
  DFFR_X1 \registers_reg[12][4]  ( .D(n3727), .CK(n675), .RN(n6785), .Q(
        \registers[12][4] ) );
  DFFR_X1 \registers_reg[12][3]  ( .D(n3726), .CK(n675), .RN(n6833), .Q(
        \registers[12][3] ) );
  DFFR_X1 \registers_reg[12][2]  ( .D(n3725), .CK(n675), .RN(n6774), .Q(
        \registers[12][2] ) );
  DFFR_X1 \registers_reg[12][1]  ( .D(n3724), .CK(n675), .RN(n6769), .Q(
        \registers[12][1] ) );
  DFFR_X1 \registers_reg[12][0]  ( .D(n3723), .CK(n675), .RN(n6855), .Q(
        \registers[12][0] ) );
  DFFR_X1 \registers_reg[13][31]  ( .D(n3722), .CK(n675), .RN(n6835), .Q(
        \registers[13][31] ) );
  DFFR_X1 \registers_reg[13][30]  ( .D(n3721), .CK(n675), .RN(n6830), .Q(
        \registers[13][30] ) );
  DFFR_X1 \registers_reg[13][29]  ( .D(n3720), .CK(n675), .RN(n6824), .Q(
        \registers[13][29] ) );
  DFFR_X1 \registers_reg[13][28]  ( .D(n3719), .CK(n675), .RN(n6819), .Q(
        \registers[13][28] ) );
  DFFR_X1 \registers_reg[13][27]  ( .D(n3718), .CK(n675), .RN(n6838), .Q(
        \registers[13][27] ) );
  DFFR_X1 \registers_reg[13][26]  ( .D(n3717), .CK(n675), .RN(n6810), .Q(
        \registers[13][26] ) );
  DFFR_X1 \registers_reg[13][25]  ( .D(n3716), .CK(n675), .RN(n6813), .Q(
        \registers[13][25] ) );
  DFFR_X1 \registers_reg[13][24]  ( .D(n3715), .CK(n675), .RN(n6805), .Q(
        \registers[13][24] ) );
  DFFR_X1 \registers_reg[13][23]  ( .D(n3714), .CK(n675), .RN(n6841), .Q(
        \registers[13][23] ) );
  DFFR_X1 \registers_reg[13][22]  ( .D(n3713), .CK(n675), .RN(n6794), .Q(
        \registers[13][22] ) );
  DFFR_X1 \registers_reg[13][21]  ( .D(n3712), .CK(n675), .RN(n6796), .Q(
        \registers[13][21] ) );
  DFFR_X1 \registers_reg[13][20]  ( .D(n3711), .CK(n675), .RN(n6788), .Q(
        \registers[13][20] ) );
  DFFR_X1 \registers_reg[13][19]  ( .D(n3710), .CK(n675), .RN(n6844), .Q(
        \registers[13][19] ) );
  DFFR_X1 \registers_reg[13][18]  ( .D(n3709), .CK(n675), .RN(n6777), .Q(
        \registers[13][18] ) );
  DFFR_X1 \registers_reg[13][17]  ( .D(n3708), .CK(n675), .RN(n6780), .Q(
        \registers[13][17] ) );
  DFFR_X1 \registers_reg[13][16]  ( .D(n3707), .CK(n675), .RN(n6771), .Q(
        \registers[13][16] ) );
  DFFR_X1 \registers_reg[13][15]  ( .D(n3706), .CK(n675), .RN(n6847), .Q(
        \registers[13][15] ) );
  DFFR_X1 \registers_reg[13][14]  ( .D(n3705), .CK(n675), .RN(n6827), .Q(
        \registers[13][14] ) );
  DFFR_X1 \registers_reg[13][13]  ( .D(n3704), .CK(n675), .RN(n6821), .Q(
        \registers[13][13] ) );
  DFFR_X1 \registers_reg[13][12]  ( .D(n3703), .CK(n675), .RN(n6816), .Q(
        \registers[13][12] ) );
  DFFR_X1 \registers_reg[13][11]  ( .D(n3702), .CK(n675), .RN(n6849), .Q(
        \registers[13][11] ) );
  DFFR_X1 \registers_reg[13][10]  ( .D(n3701), .CK(n675), .RN(n6808), .Q(
        \registers[13][10] ) );
  DFFR_X1 \registers_reg[13][9]  ( .D(n3700), .CK(n675), .RN(n6799), .Q(
        \registers[13][9] ) );
  DFFR_X1 \registers_reg[13][8]  ( .D(n3699), .CK(n675), .RN(n6802), .Q(
        \registers[13][8] ) );
  DFFR_X1 \registers_reg[13][7]  ( .D(n3698), .CK(n675), .RN(n6852), .Q(
        \registers[13][7] ) );
  DFFR_X1 \registers_reg[13][6]  ( .D(n3697), .CK(n675), .RN(n6791), .Q(
        \registers[13][6] ) );
  DFFR_X1 \registers_reg[13][5]  ( .D(n3696), .CK(n675), .RN(n6783), .Q(
        \registers[13][5] ) );
  DFFR_X1 \registers_reg[13][4]  ( .D(n3695), .CK(n675), .RN(n6785), .Q(
        \registers[13][4] ) );
  DFFR_X1 \registers_reg[13][3]  ( .D(n3694), .CK(n675), .RN(n6832), .Q(
        \registers[13][3] ) );
  DFFR_X1 \registers_reg[13][2]  ( .D(n3693), .CK(n675), .RN(n6774), .Q(
        \registers[13][2] ) );
  DFFR_X1 \registers_reg[13][1]  ( .D(n3692), .CK(n675), .RN(n6769), .Q(
        \registers[13][1] ) );
  DFFR_X1 \registers_reg[13][0]  ( .D(n3691), .CK(n675), .RN(n6855), .Q(
        \registers[13][0] ) );
  DFFR_X1 \registers_reg[14][31]  ( .D(n3690), .CK(n675), .RN(n6835), .Q(
        \registers[14][31] ) );
  DFFR_X1 \registers_reg[14][30]  ( .D(n3689), .CK(n675), .RN(n6830), .Q(
        \registers[14][30] ) );
  DFFR_X1 \registers_reg[14][29]  ( .D(n3688), .CK(n675), .RN(n6824), .Q(
        \registers[14][29] ) );
  DFFR_X1 \registers_reg[14][28]  ( .D(n3687), .CK(n675), .RN(n6819), .Q(
        \registers[14][28] ) );
  DFFR_X1 \registers_reg[14][27]  ( .D(n3686), .CK(n675), .RN(n6838), .Q(
        \registers[14][27] ) );
  DFFR_X1 \registers_reg[14][26]  ( .D(n3685), .CK(n675), .RN(n6810), .Q(
        \registers[14][26] ) );
  DFFR_X1 \registers_reg[14][25]  ( .D(n3684), .CK(n675), .RN(n6813), .Q(
        \registers[14][25] ) );
  DFFR_X1 \registers_reg[14][24]  ( .D(n3683), .CK(n675), .RN(n6805), .Q(
        \registers[14][24] ) );
  DFFR_X1 \registers_reg[14][23]  ( .D(n3682), .CK(n675), .RN(n6841), .Q(
        \registers[14][23] ) );
  DFFR_X1 \registers_reg[14][22]  ( .D(n3681), .CK(n675), .RN(n6794), .Q(
        \registers[14][22] ) );
  DFFR_X1 \registers_reg[14][21]  ( .D(n3680), .CK(n675), .RN(n6796), .Q(
        \registers[14][21] ) );
  DFFR_X1 \registers_reg[14][20]  ( .D(n3679), .CK(n675), .RN(n6788), .Q(
        \registers[14][20] ) );
  DFFR_X1 \registers_reg[14][19]  ( .D(n3678), .CK(n675), .RN(n6844), .Q(
        \registers[14][19] ) );
  DFFR_X1 \registers_reg[14][18]  ( .D(n3677), .CK(n675), .RN(n6777), .Q(
        \registers[14][18] ) );
  DFFR_X1 \registers_reg[14][17]  ( .D(n3676), .CK(n675), .RN(n6780), .Q(
        \registers[14][17] ) );
  DFFR_X1 \registers_reg[14][16]  ( .D(n3675), .CK(n675), .RN(n6771), .Q(
        \registers[14][16] ) );
  DFFR_X1 \registers_reg[14][15]  ( .D(n3674), .CK(n675), .RN(n6846), .Q(
        \registers[14][15] ) );
  DFFR_X1 \registers_reg[14][14]  ( .D(n3673), .CK(n675), .RN(n6827), .Q(
        \registers[14][14] ) );
  DFFR_X1 \registers_reg[14][13]  ( .D(n3672), .CK(n675), .RN(n6821), .Q(
        \registers[14][13] ) );
  DFFR_X1 \registers_reg[14][12]  ( .D(n3671), .CK(n675), .RN(n6816), .Q(
        \registers[14][12] ) );
  DFFR_X1 \registers_reg[14][11]  ( .D(n3670), .CK(n675), .RN(n6849), .Q(
        \registers[14][11] ) );
  DFFR_X1 \registers_reg[14][10]  ( .D(n3669), .CK(n675), .RN(n6807), .Q(
        \registers[14][10] ) );
  DFFR_X1 \registers_reg[14][9]  ( .D(n3668), .CK(n675), .RN(n6799), .Q(
        \registers[14][9] ) );
  DFFR_X1 \registers_reg[14][8]  ( .D(n3667), .CK(n675), .RN(n6802), .Q(
        \registers[14][8] ) );
  DFFR_X1 \registers_reg[14][7]  ( .D(n3666), .CK(n675), .RN(n6852), .Q(
        \registers[14][7] ) );
  DFFR_X1 \registers_reg[14][6]  ( .D(n3665), .CK(n675), .RN(n6791), .Q(
        \registers[14][6] ) );
  DFFR_X1 \registers_reg[14][5]  ( .D(n3664), .CK(n675), .RN(n6782), .Q(
        \registers[14][5] ) );
  DFFR_X1 \registers_reg[14][4]  ( .D(n3663), .CK(n675), .RN(n6785), .Q(
        \registers[14][4] ) );
  DFFR_X1 \registers_reg[14][3]  ( .D(n3662), .CK(n675), .RN(n6832), .Q(
        \registers[14][3] ) );
  DFFR_X1 \registers_reg[14][2]  ( .D(n3661), .CK(n675), .RN(n6774), .Q(
        \registers[14][2] ) );
  DFFR_X1 \registers_reg[14][1]  ( .D(n3660), .CK(n675), .RN(n6769), .Q(
        \registers[14][1] ) );
  DFFR_X1 \registers_reg[14][0]  ( .D(n3659), .CK(n675), .RN(n6855), .Q(
        \registers[14][0] ) );
  DFFR_X1 \registers_reg[15][31]  ( .D(n3658), .CK(n675), .RN(n6835), .Q(
        \registers[15][31] ) );
  DFFR_X1 \registers_reg[15][30]  ( .D(n3657), .CK(n675), .RN(n6829), .Q(
        \registers[15][30] ) );
  DFFR_X1 \registers_reg[15][29]  ( .D(n3656), .CK(n675), .RN(n6824), .Q(
        \registers[15][29] ) );
  DFFR_X1 \registers_reg[15][28]  ( .D(n3655), .CK(n675), .RN(n6818), .Q(
        \registers[15][28] ) );
  DFFR_X1 \registers_reg[15][27]  ( .D(n3654), .CK(n675), .RN(n6838), .Q(
        \registers[15][27] ) );
  DFFR_X1 \registers_reg[15][26]  ( .D(n3653), .CK(n675), .RN(n6810), .Q(
        \registers[15][26] ) );
  DFFR_X1 \registers_reg[15][25]  ( .D(n3652), .CK(n675), .RN(n6813), .Q(
        \registers[15][25] ) );
  DFFR_X1 \registers_reg[15][24]  ( .D(n3651), .CK(n675), .RN(n6805), .Q(
        \registers[15][24] ) );
  DFFR_X1 \registers_reg[15][23]  ( .D(n3650), .CK(n675), .RN(n6841), .Q(
        \registers[15][23] ) );
  DFFR_X1 \registers_reg[15][22]  ( .D(n3649), .CK(n675), .RN(n6793), .Q(
        \registers[15][22] ) );
  DFFR_X1 \registers_reg[15][21]  ( .D(n3648), .CK(n675), .RN(n6796), .Q(
        \registers[15][21] ) );
  DFFR_X1 \registers_reg[15][20]  ( .D(n3647), .CK(n675), .RN(n6788), .Q(
        \registers[15][20] ) );
  DFFR_X1 \registers_reg[15][19]  ( .D(n3646), .CK(n675), .RN(n6844), .Q(
        \registers[15][19] ) );
  DFFR_X1 \registers_reg[15][18]  ( .D(n3645), .CK(n675), .RN(n6777), .Q(
        \registers[15][18] ) );
  DFFR_X1 \registers_reg[15][17]  ( .D(n3644), .CK(n675), .RN(n6780), .Q(
        \registers[15][17] ) );
  DFFR_X1 \registers_reg[15][16]  ( .D(n3643), .CK(n675), .RN(n6771), .Q(
        \registers[15][16] ) );
  DFFR_X1 \registers_reg[15][15]  ( .D(n3642), .CK(n675), .RN(n6846), .Q(
        \registers[15][15] ) );
  DFFR_X1 \registers_reg[15][14]  ( .D(n3641), .CK(n675), .RN(n6827), .Q(
        \registers[15][14] ) );
  DFFR_X1 \registers_reg[15][13]  ( .D(n3640), .CK(n675), .RN(n6821), .Q(
        \registers[15][13] ) );
  DFFR_X1 \registers_reg[15][12]  ( .D(n3639), .CK(n675), .RN(n6816), .Q(
        \registers[15][12] ) );
  DFFR_X1 \registers_reg[15][11]  ( .D(n3638), .CK(n675), .RN(n6849), .Q(
        \registers[15][11] ) );
  DFFR_X1 \registers_reg[15][10]  ( .D(n3637), .CK(n675), .RN(n6807), .Q(
        \registers[15][10] ) );
  DFFR_X1 \registers_reg[15][9]  ( .D(n3636), .CK(n675), .RN(n6799), .Q(
        \registers[15][9] ) );
  DFFR_X1 \registers_reg[15][8]  ( .D(n3635), .CK(n675), .RN(n6802), .Q(
        \registers[15][8] ) );
  DFFR_X1 \registers_reg[15][7]  ( .D(n3634), .CK(n675), .RN(n6852), .Q(
        \registers[15][7] ) );
  DFFR_X1 \registers_reg[15][6]  ( .D(n3633), .CK(n675), .RN(n6791), .Q(
        \registers[15][6] ) );
  DFFR_X1 \registers_reg[15][5]  ( .D(n3632), .CK(n675), .RN(n6782), .Q(
        \registers[15][5] ) );
  DFFR_X1 \registers_reg[15][4]  ( .D(n3631), .CK(n675), .RN(n6785), .Q(
        \registers[15][4] ) );
  DFFR_X1 \registers_reg[15][3]  ( .D(n3630), .CK(n675), .RN(n6832), .Q(
        \registers[15][3] ) );
  DFFR_X1 \registers_reg[15][2]  ( .D(n3629), .CK(n675), .RN(n6774), .Q(
        \registers[15][2] ) );
  DFFR_X1 \registers_reg[15][1]  ( .D(n3628), .CK(n675), .RN(n6768), .Q(
        \registers[15][1] ) );
  DFFR_X1 \registers_reg[15][0]  ( .D(n3627), .CK(n675), .RN(n6855), .Q(
        \registers[15][0] ) );
  DFFR_X1 \registers_reg[16][31]  ( .D(n3626), .CK(n675), .RN(n6835), .Q(
        \registers[16][31] ), .QN(n5841) );
  DFFR_X1 \registers_reg[16][30]  ( .D(n3625), .CK(n675), .RN(n6829), .Q(
        \registers[16][30] ), .QN(n5839) );
  DFFR_X1 \registers_reg[16][29]  ( .D(n3624), .CK(n675), .RN(n6824), .Q(
        \registers[16][29] ), .QN(n5837) );
  DFFR_X1 \registers_reg[16][28]  ( .D(n3623), .CK(n675), .RN(n6818), .Q(
        \registers[16][28] ), .QN(n5835) );
  DFFR_X1 \registers_reg[16][27]  ( .D(n3622), .CK(n675), .RN(n6838), .Q(
        \registers[16][27] ), .QN(n5917) );
  DFFR_X1 \registers_reg[16][26]  ( .D(n3621), .CK(n675), .RN(n6810), .Q(
        \registers[16][26] ), .QN(n5916) );
  DFFR_X1 \registers_reg[16][25]  ( .D(n3620), .CK(n675), .RN(n6813), .Q(
        \registers[16][25] ), .QN(n5915) );
  DFFR_X1 \registers_reg[16][24]  ( .D(n3619), .CK(n675), .RN(n6805), .Q(
        \registers[16][24] ), .QN(n5914) );
  DFFR_X1 \registers_reg[16][23]  ( .D(n3618), .CK(n675), .RN(n6841), .Q(
        \registers[16][23] ), .QN(n5913) );
  DFFR_X1 \registers_reg[16][22]  ( .D(n3617), .CK(n675), .RN(n6793), .Q(
        \registers[16][22] ), .QN(n5912) );
  DFFR_X1 \registers_reg[16][21]  ( .D(n3616), .CK(n675), .RN(n6796), .Q(
        \registers[16][21] ), .QN(n5827) );
  DFFR_X1 \registers_reg[16][20]  ( .D(n3615), .CK(n675), .RN(n6788), .Q(
        \registers[16][20] ), .QN(n5825) );
  DFFR_X1 \registers_reg[16][19]  ( .D(n3614), .CK(n675), .RN(n6843), .Q(
        \registers[16][19] ), .QN(n5823) );
  DFFR_X1 \registers_reg[16][18]  ( .D(n3613), .CK(n675), .RN(n6777), .Q(
        \registers[16][18] ), .QN(n5821) );
  DFFR_X1 \registers_reg[16][17]  ( .D(n3612), .CK(n675), .RN(n6780), .Q(
        \registers[16][17] ), .QN(n5819) );
  DFFR_X1 \registers_reg[16][16]  ( .D(n3611), .CK(n675), .RN(n6771), .Q(
        \registers[16][16] ), .QN(n5817) );
  DFFR_X1 \registers_reg[16][15]  ( .D(n3610), .CK(n675), .RN(n6846), .Q(
        \registers[16][15] ), .QN(n5815) );
  DFFR_X1 \registers_reg[16][14]  ( .D(n3609), .CK(n675), .RN(n6827), .Q(
        \registers[16][14] ), .QN(n5813) );
  DFFR_X1 \registers_reg[16][13]  ( .D(n3608), .CK(n675), .RN(n6821), .Q(
        \registers[16][13] ), .QN(n5811) );
  DFFR_X1 \registers_reg[16][12]  ( .D(n3607), .CK(n675), .RN(n6816), .Q(
        \registers[16][12] ), .QN(n5809) );
  DFFR_X1 \registers_reg[16][11]  ( .D(n3606), .CK(n675), .RN(n6849), .Q(
        \registers[16][11] ), .QN(n5807) );
  DFFR_X1 \registers_reg[16][10]  ( .D(n3605), .CK(n675), .RN(n6807), .Q(
        \registers[16][10] ), .QN(n5805) );
  DFFR_X1 \registers_reg[16][9]  ( .D(n3604), .CK(n675), .RN(n6799), .Q(
        \registers[16][9] ), .QN(n5803) );
  DFFR_X1 \registers_reg[16][8]  ( .D(n3603), .CK(n675), .RN(n6802), .Q(
        \registers[16][8] ), .QN(n5801) );
  DFFR_X1 \registers_reg[16][7]  ( .D(n3602), .CK(n675), .RN(n6852), .Q(
        \registers[16][7] ), .QN(n5799) );
  DFFR_X1 \registers_reg[16][6]  ( .D(n3601), .CK(n675), .RN(n6791), .Q(
        \registers[16][6] ), .QN(n5797) );
  DFFR_X1 \registers_reg[16][5]  ( .D(n3600), .CK(n675), .RN(n6782), .Q(
        \registers[16][5] ), .QN(n5795) );
  DFFR_X1 \registers_reg[16][4]  ( .D(n3599), .CK(n675), .RN(n6785), .Q(
        \registers[16][4] ), .QN(n5793) );
  DFFR_X1 \registers_reg[16][3]  ( .D(n3598), .CK(n675), .RN(n6832), .Q(
        \registers[16][3] ), .QN(n5791) );
  DFFR_X1 \registers_reg[16][2]  ( .D(n3597), .CK(n675), .RN(n6774), .Q(
        \registers[16][2] ), .QN(n5789) );
  DFFR_X1 \registers_reg[16][1]  ( .D(n3596), .CK(n675), .RN(n6768), .Q(
        \registers[16][1] ), .QN(n5787) );
  DFFR_X1 \registers_reg[16][0]  ( .D(n3595), .CK(n675), .RN(n6855), .Q(
        \registers[16][0] ), .QN(n5785) );
  DFFR_X1 \registers_reg[17][31]  ( .D(n3594), .CK(n675), .RN(n6835), .Q(
        \registers[17][31] ), .QN(n2851) );
  DFFR_X1 \registers_reg[17][30]  ( .D(n3593), .CK(n675), .RN(n6829), .Q(
        \registers[17][30] ), .QN(n2849) );
  DFFR_X1 \registers_reg[17][29]  ( .D(n3592), .CK(n675), .RN(n6824), .Q(
        \registers[17][29] ), .QN(n2847) );
  DFFR_X1 \registers_reg[17][28]  ( .D(n3591), .CK(n675), .RN(n6818), .Q(
        \registers[17][28] ), .QN(n2845) );
  DFFR_X1 \registers_reg[17][27]  ( .D(n3590), .CK(n675), .RN(n6838), .Q(
        \registers[17][27] ), .QN(n4219) );
  DFFR_X1 \registers_reg[17][26]  ( .D(n3589), .CK(n675), .RN(n6810), .Q(
        \registers[17][26] ), .QN(n4218) );
  DFFR_X1 \registers_reg[17][25]  ( .D(n3588), .CK(n675), .RN(n6813), .Q(
        \registers[17][25] ), .QN(n4216) );
  DFFR_X1 \registers_reg[17][24]  ( .D(n3587), .CK(n675), .RN(n6804), .Q(
        \registers[17][24] ), .QN(n4215) );
  DFFR_X1 \registers_reg[17][23]  ( .D(n3586), .CK(n675), .RN(n6841), .Q(
        \registers[17][23] ), .QN(n4214) );
  DFFR_X1 \registers_reg[17][22]  ( .D(n3585), .CK(n675), .RN(n6793), .Q(
        \registers[17][22] ), .QN(n4213) );
  DFFR_X1 \registers_reg[17][21]  ( .D(n3584), .CK(n675), .RN(n6796), .Q(
        \registers[17][21] ), .QN(n2837) );
  DFFR_X1 \registers_reg[17][20]  ( .D(n3583), .CK(n675), .RN(n6788), .Q(
        \registers[17][20] ), .QN(n2835) );
  DFFR_X1 \registers_reg[17][19]  ( .D(n3582), .CK(n675), .RN(n6843), .Q(
        \registers[17][19] ), .QN(n2833) );
  DFFR_X1 \registers_reg[17][18]  ( .D(n3581), .CK(n675), .RN(n6777), .Q(
        \registers[17][18] ), .QN(n2831) );
  DFFR_X1 \registers_reg[17][17]  ( .D(n3580), .CK(n675), .RN(n6779), .Q(
        \registers[17][17] ), .QN(n2829) );
  DFFR_X1 \registers_reg[17][16]  ( .D(n3579), .CK(n675), .RN(n6771), .Q(
        \registers[17][16] ), .QN(n2827) );
  DFFR_X1 \registers_reg[17][15]  ( .D(n3578), .CK(n675), .RN(n6846), .Q(
        \registers[17][15] ), .QN(n2823) );
  DFFR_X1 \registers_reg[17][14]  ( .D(n3577), .CK(n675), .RN(n6827), .Q(
        \registers[17][14] ), .QN(n2821) );
  DFFR_X1 \registers_reg[17][13]  ( .D(n3576), .CK(n675), .RN(n6821), .Q(
        \registers[17][13] ), .QN(n2819) );
  DFFR_X1 \registers_reg[17][12]  ( .D(n3575), .CK(n675), .RN(n6816), .Q(
        \registers[17][12] ), .QN(n2817) );
  DFFR_X1 \registers_reg[17][11]  ( .D(n3574), .CK(n675), .RN(n6849), .Q(
        \registers[17][11] ), .QN(n2815) );
  DFFR_X1 \registers_reg[17][10]  ( .D(n3573), .CK(n675), .RN(n6807), .Q(
        \registers[17][10] ), .QN(n2813) );
  DFFR_X1 \registers_reg[17][9]  ( .D(n3572), .CK(n675), .RN(n6799), .Q(
        \registers[17][9] ), .QN(n2811) );
  DFFR_X1 \registers_reg[17][8]  ( .D(n3571), .CK(n675), .RN(n6802), .Q(
        \registers[17][8] ), .QN(n2809) );
  DFFR_X1 \registers_reg[17][7]  ( .D(n3570), .CK(n675), .RN(n6852), .Q(
        \registers[17][7] ), .QN(n2807) );
  DFFR_X1 \registers_reg[17][6]  ( .D(n3569), .CK(n675), .RN(n6791), .Q(
        \registers[17][6] ), .QN(n2805) );
  DFFR_X1 \registers_reg[17][5]  ( .D(n3568), .CK(n675), .RN(n6782), .Q(
        \registers[17][5] ), .QN(n2803) );
  DFFR_X1 \registers_reg[17][4]  ( .D(n3567), .CK(n675), .RN(n6785), .Q(
        \registers[17][4] ), .QN(n2801) );
  DFFR_X1 \registers_reg[17][3]  ( .D(n3566), .CK(n675), .RN(n6832), .Q(
        \registers[17][3] ), .QN(n2799) );
  DFFR_X1 \registers_reg[17][2]  ( .D(n3565), .CK(n675), .RN(n6774), .Q(
        \registers[17][2] ), .QN(n2797) );
  DFFR_X1 \registers_reg[17][1]  ( .D(n3564), .CK(n675), .RN(n6768), .Q(
        \registers[17][1] ), .QN(n2795) );
  DFFR_X1 \registers_reg[17][0]  ( .D(n3563), .CK(n675), .RN(n6855), .Q(
        \registers[17][0] ), .QN(n2793) );
  DFFR_X1 \registers_reg[18][31]  ( .D(n3562), .CK(n675), .RN(n6835), .Q(
        \registers[18][31] ), .QN(n5897) );
  DFFR_X1 \registers_reg[18][30]  ( .D(n3561), .CK(n675), .RN(n6829), .Q(
        \registers[18][30] ), .QN(n5895) );
  DFFR_X1 \registers_reg[18][29]  ( .D(n3560), .CK(n675), .RN(n6824), .Q(
        \registers[18][29] ), .QN(n5893) );
  DFFR_X1 \registers_reg[18][28]  ( .D(n3559), .CK(n675), .RN(n6818), .Q(
        \registers[18][28] ), .QN(n5891) );
  DFFR_X1 \registers_reg[18][27]  ( .D(n3558), .CK(n675), .RN(n6838), .Q(
        \registers[18][27] ), .QN(n5889) );
  DFFR_X1 \registers_reg[18][26]  ( .D(n3557), .CK(n675), .RN(n6810), .Q(
        \registers[18][26] ), .QN(n5888) );
  DFFR_X1 \registers_reg[18][25]  ( .D(n3556), .CK(n675), .RN(n6813), .Q(
        \registers[18][25] ), .QN(n5887) );
  DFFR_X1 \registers_reg[18][24]  ( .D(n3555), .CK(n675), .RN(n6804), .Q(
        \registers[18][24] ), .QN(n5886) );
  DFFR_X1 \registers_reg[18][23]  ( .D(n3554), .CK(n675), .RN(n6840), .Q(
        \registers[18][23] ), .QN(n5885) );
  DFFR_X1 \registers_reg[18][22]  ( .D(n3553), .CK(n675), .RN(n6793), .Q(
        \registers[18][22] ), .QN(n5884) );
  DFFR_X1 \registers_reg[18][21]  ( .D(n3552), .CK(n675), .RN(n6796), .Q(
        \registers[18][21] ), .QN(n5883) );
  DFFR_X1 \registers_reg[18][20]  ( .D(n3551), .CK(n675), .RN(n6788), .Q(
        \registers[18][20] ), .QN(n5882) );
  DFFR_X1 \registers_reg[18][19]  ( .D(n3550), .CK(n675), .RN(n6843), .Q(
        \registers[18][19] ), .QN(n5881) );
  DFFR_X1 \registers_reg[18][18]  ( .D(n3549), .CK(n675), .RN(n6777), .Q(
        \registers[18][18] ), .QN(n5879) );
  DFFR_X1 \registers_reg[18][17]  ( .D(n3548), .CK(n675), .RN(n6779), .Q(
        \registers[18][17] ), .QN(n5877) );
  DFFR_X1 \registers_reg[18][16]  ( .D(n3547), .CK(n675), .RN(n6771), .Q(
        \registers[18][16] ), .QN(n5875) );
  DFFR_X1 \registers_reg[18][15]  ( .D(n3546), .CK(n675), .RN(n6846), .Q(
        \registers[18][15] ), .QN(n5873) );
  DFFR_X1 \registers_reg[18][14]  ( .D(n3545), .CK(n675), .RN(n6826), .Q(
        \registers[18][14] ), .QN(n5871) );
  DFFR_X1 \registers_reg[18][13]  ( .D(n3544), .CK(n675), .RN(n6821), .Q(
        \registers[18][13] ), .QN(n5869) );
  DFFR_X1 \registers_reg[18][12]  ( .D(n3543), .CK(n675), .RN(n6815), .Q(
        \registers[18][12] ), .QN(n5867) );
  DFFR_X1 \registers_reg[18][11]  ( .D(n3542), .CK(n675), .RN(n6849), .Q(
        \registers[18][11] ), .QN(n5865) );
  DFFR_X1 \registers_reg[18][10]  ( .D(n3541), .CK(n675), .RN(n6807), .Q(
        \registers[18][10] ), .QN(n5863) );
  DFFR_X1 \registers_reg[18][9]  ( .D(n3540), .CK(n675), .RN(n6799), .Q(
        \registers[18][9] ), .QN(n5861) );
  DFFR_X1 \registers_reg[18][8]  ( .D(n3539), .CK(n675), .RN(n6802), .Q(
        \registers[18][8] ), .QN(n5859) );
  DFFR_X1 \registers_reg[18][7]  ( .D(n3538), .CK(n675), .RN(n6852), .Q(
        \registers[18][7] ), .QN(n5857) );
  DFFR_X1 \registers_reg[18][6]  ( .D(n3537), .CK(n675), .RN(n6790), .Q(
        \registers[18][6] ), .QN(n5855) );
  DFFR_X1 \registers_reg[18][5]  ( .D(n3536), .CK(n675), .RN(n6782), .Q(
        \registers[18][5] ), .QN(n5853) );
  DFFR_X1 \registers_reg[18][4]  ( .D(n3535), .CK(n675), .RN(n6785), .Q(
        \registers[18][4] ), .QN(n5851) );
  DFFR_X1 \registers_reg[18][3]  ( .D(n3534), .CK(n675), .RN(n6832), .Q(
        \registers[18][3] ), .QN(n5849) );
  DFFR_X1 \registers_reg[18][2]  ( .D(n3533), .CK(n675), .RN(n6774), .Q(
        \registers[18][2] ), .QN(n5847) );
  DFFR_X1 \registers_reg[18][1]  ( .D(n3532), .CK(n675), .RN(n6768), .Q(
        \registers[18][1] ), .QN(n5845) );
  DFFR_X1 \registers_reg[18][0]  ( .D(n3531), .CK(n675), .RN(n6855), .Q(
        \registers[18][0] ), .QN(n5843) );
  DFFR_X1 \registers_reg[19][31]  ( .D(n3530), .CK(n675), .RN(n6835), .Q(
        \registers[19][31] ), .QN(n4198) );
  DFFR_X1 \registers_reg[19][30]  ( .D(n3529), .CK(n675), .RN(n6829), .Q(
        \registers[19][30] ), .QN(n4196) );
  DFFR_X1 \registers_reg[19][29]  ( .D(n3528), .CK(n675), .RN(n6824), .Q(
        \registers[19][29] ), .QN(n4194) );
  DFFR_X1 \registers_reg[19][28]  ( .D(n3527), .CK(n675), .RN(n6818), .Q(
        \registers[19][28] ), .QN(n4192) );
  DFFR_X1 \registers_reg[19][27]  ( .D(n3526), .CK(n675), .RN(n6838), .Q(
        \registers[19][27] ), .QN(n4190) );
  DFFR_X1 \registers_reg[19][26]  ( .D(n3525), .CK(n675), .RN(n6810), .Q(
        \registers[19][26] ), .QN(n4189) );
  DFFR_X1 \registers_reg[19][25]  ( .D(n3524), .CK(n675), .RN(n6813), .Q(
        \registers[19][25] ), .QN(n4188) );
  DFFR_X1 \registers_reg[19][24]  ( .D(n3523), .CK(n675), .RN(n6804), .Q(
        \registers[19][24] ), .QN(n4187) );
  DFFR_X1 \registers_reg[19][23]  ( .D(n3522), .CK(n675), .RN(n6840), .Q(
        \registers[19][23] ), .QN(n4186) );
  DFFR_X1 \registers_reg[19][22]  ( .D(n3521), .CK(n675), .RN(n6793), .Q(
        \registers[19][22] ), .QN(n4185) );
  DFFR_X1 \registers_reg[19][21]  ( .D(n3520), .CK(n675), .RN(n6796), .Q(
        \registers[19][21] ), .QN(n4181) );
  DFFR_X1 \registers_reg[19][20]  ( .D(n3519), .CK(n675), .RN(n6788), .Q(
        \registers[19][20] ), .QN(n4180) );
  DFFR_X1 \registers_reg[19][19]  ( .D(n3518), .CK(n675), .RN(n6843), .Q(
        \registers[19][19] ), .QN(n4179) );
  DFFR_X1 \registers_reg[19][18]  ( .D(n3517), .CK(n675), .RN(n6776), .Q(
        \registers[19][18] ), .QN(n4177) );
  DFFR_X1 \registers_reg[19][17]  ( .D(n3516), .CK(n675), .RN(n6779), .Q(
        \registers[19][17] ), .QN(n4175) );
  DFFR_X1 \registers_reg[19][16]  ( .D(n3515), .CK(n675), .RN(n6771), .Q(
        \registers[19][16] ), .QN(n4173) );
  DFFR_X1 \registers_reg[19][15]  ( .D(n3514), .CK(n675), .RN(n6846), .Q(
        \registers[19][15] ), .QN(n4171) );
  DFFR_X1 \registers_reg[19][14]  ( .D(n3513), .CK(n675), .RN(n6826), .Q(
        \registers[19][14] ), .QN(n4169) );
  DFFR_X1 \registers_reg[19][13]  ( .D(n3512), .CK(n675), .RN(n6821), .Q(
        \registers[19][13] ), .QN(n4167) );
  DFFR_X1 \registers_reg[19][12]  ( .D(n3511), .CK(n675), .RN(n6815), .Q(
        \registers[19][12] ), .QN(n4165) );
  DFFR_X1 \registers_reg[19][11]  ( .D(n3510), .CK(n675), .RN(n6849), .Q(
        \registers[19][11] ), .QN(n4163) );
  DFFR_X1 \registers_reg[19][10]  ( .D(n3509), .CK(n675), .RN(n6807), .Q(
        \registers[19][10] ), .QN(n4161) );
  DFFR_X1 \registers_reg[19][9]  ( .D(n3508), .CK(n675), .RN(n6799), .Q(
        \registers[19][9] ), .QN(n4159) );
  DFFR_X1 \registers_reg[19][8]  ( .D(n3507), .CK(n675), .RN(n6802), .Q(
        \registers[19][8] ), .QN(n4157) );
  DFFR_X1 \registers_reg[19][7]  ( .D(n3506), .CK(n675), .RN(n6852), .Q(
        \registers[19][7] ), .QN(n4155) );
  DFFR_X1 \registers_reg[19][6]  ( .D(n3505), .CK(n675), .RN(n6790), .Q(
        \registers[19][6] ), .QN(n4153) );
  DFFR_X1 \registers_reg[19][5]  ( .D(n3504), .CK(n675), .RN(n6782), .Q(
        \registers[19][5] ), .QN(n4151) );
  DFFR_X1 \registers_reg[19][4]  ( .D(n3503), .CK(n675), .RN(n6785), .Q(
        \registers[19][4] ), .QN(n2971) );
  DFFR_X1 \registers_reg[19][3]  ( .D(n3502), .CK(n675), .RN(n6832), .Q(
        \registers[19][3] ), .QN(n2895) );
  DFFR_X1 \registers_reg[19][2]  ( .D(n3501), .CK(n675), .RN(n6774), .Q(
        \registers[19][2] ), .QN(n2857) );
  DFFR_X1 \registers_reg[19][1]  ( .D(n3500), .CK(n675), .RN(n6768), .Q(
        \registers[19][1] ), .QN(n2855) );
  DFFR_X1 \registers_reg[19][0]  ( .D(n3499), .CK(n675), .RN(n6855), .Q(
        \registers[19][0] ), .QN(n2853) );
  DFFR_X1 \registers_reg[20][31]  ( .D(n3498), .CK(n675), .RN(n6835), .Q(
        \registers[20][31] ) );
  DFFR_X1 \registers_reg[20][30]  ( .D(n3497), .CK(n675), .RN(n6829), .Q(
        \registers[20][30] ) );
  DFFR_X1 \registers_reg[20][29]  ( .D(n3496), .CK(n675), .RN(n6824), .Q(
        \registers[20][29] ) );
  DFFR_X1 \registers_reg[20][28]  ( .D(n3495), .CK(n675), .RN(n6818), .Q(
        \registers[20][28] ) );
  DFFR_X1 \registers_reg[20][27]  ( .D(n3494), .CK(n675), .RN(n6837), .Q(
        \registers[20][27] ) );
  DFFR_X1 \registers_reg[20][26]  ( .D(n3493), .CK(n675), .RN(n6810), .Q(
        \registers[20][26] ) );
  DFFR_X1 \registers_reg[20][25]  ( .D(n3492), .CK(n675), .RN(n6813), .Q(
        \registers[20][25] ) );
  DFFR_X1 \registers_reg[20][24]  ( .D(n3491), .CK(n675), .RN(n6804), .Q(
        \registers[20][24] ) );
  DFFR_X1 \registers_reg[20][23]  ( .D(n3490), .CK(n675), .RN(n6840), .Q(
        \registers[20][23] ) );
  DFFR_X1 \registers_reg[20][22]  ( .D(n3489), .CK(n675), .RN(n6793), .Q(
        \registers[20][22] ) );
  DFFR_X1 \registers_reg[20][21]  ( .D(n3488), .CK(n675), .RN(n6796), .Q(
        \registers[20][21] ) );
  DFFR_X1 \registers_reg[20][20]  ( .D(n3487), .CK(n675), .RN(n6788), .Q(
        \registers[20][20] ) );
  DFFR_X1 \registers_reg[20][19]  ( .D(n3486), .CK(n675), .RN(n6843), .Q(
        \registers[20][19] ) );
  DFFR_X1 \registers_reg[20][18]  ( .D(n3485), .CK(n675), .RN(n6776), .Q(
        \registers[20][18] ) );
  DFFR_X1 \registers_reg[20][17]  ( .D(n3484), .CK(n675), .RN(n6779), .Q(
        \registers[20][17] ) );
  DFFR_X1 \registers_reg[20][16]  ( .D(n3483), .CK(n675), .RN(n6771), .Q(
        \registers[20][16] ) );
  DFFR_X1 \registers_reg[20][15]  ( .D(n3482), .CK(n675), .RN(n6846), .Q(
        \registers[20][15] ) );
  DFFR_X1 \registers_reg[20][14]  ( .D(n3481), .CK(n675), .RN(n6826), .Q(
        \registers[20][14] ) );
  DFFR_X1 \registers_reg[20][13]  ( .D(n3480), .CK(n675), .RN(n6821), .Q(
        \registers[20][13] ) );
  DFFR_X1 \registers_reg[20][12]  ( .D(n3479), .CK(n675), .RN(n6815), .Q(
        \registers[20][12] ) );
  DFFR_X1 \registers_reg[20][11]  ( .D(n3478), .CK(n675), .RN(n6849), .Q(
        \registers[20][11] ) );
  DFFR_X1 \registers_reg[20][10]  ( .D(n3477), .CK(n675), .RN(n6807), .Q(
        \registers[20][10] ) );
  DFFR_X1 \registers_reg[20][9]  ( .D(n3476), .CK(n675), .RN(n6799), .Q(
        \registers[20][9] ) );
  DFFR_X1 \registers_reg[20][8]  ( .D(n3475), .CK(n675), .RN(n6801), .Q(
        \registers[20][8] ) );
  DFFR_X1 \registers_reg[20][7]  ( .D(n3474), .CK(n675), .RN(n6852), .Q(
        \registers[20][7] ) );
  DFFR_X1 \registers_reg[20][6]  ( .D(n3473), .CK(n675), .RN(n6790), .Q(
        \registers[20][6] ) );
  DFFR_X1 \registers_reg[20][5]  ( .D(n3472), .CK(n675), .RN(n6782), .Q(
        \registers[20][5] ) );
  DFFR_X1 \registers_reg[20][4]  ( .D(n3471), .CK(n675), .RN(n6785), .Q(
        \registers[20][4] ) );
  DFFR_X1 \registers_reg[20][3]  ( .D(n3470), .CK(n675), .RN(n6832), .Q(
        \registers[20][3] ) );
  DFFR_X1 \registers_reg[20][2]  ( .D(n3469), .CK(n675), .RN(n6774), .Q(
        \registers[20][2] ) );
  DFFR_X1 \registers_reg[20][1]  ( .D(n3468), .CK(n675), .RN(n6768), .Q(
        \registers[20][1] ) );
  DFFR_X1 \registers_reg[20][0]  ( .D(n3467), .CK(n675), .RN(n6854), .Q(
        \registers[20][0] ) );
  DFFR_X1 \registers_reg[21][31]  ( .D(n3466), .CK(n675), .RN(n6835), .Q(
        \registers[21][31] ) );
  DFFR_X1 \registers_reg[21][30]  ( .D(n3465), .CK(n675), .RN(n6829), .Q(
        \registers[21][30] ) );
  DFFR_X1 \registers_reg[21][29]  ( .D(n3464), .CK(n675), .RN(n6823), .Q(
        \registers[21][29] ) );
  DFFR_X1 \registers_reg[21][28]  ( .D(n3463), .CK(n675), .RN(n6818), .Q(
        \registers[21][28] ) );
  DFFR_X1 \registers_reg[21][27]  ( .D(n3462), .CK(n675), .RN(n6837), .Q(
        \registers[21][27] ) );
  DFFR_X1 \registers_reg[21][26]  ( .D(n3461), .CK(n675), .RN(n6810), .Q(
        \registers[21][26] ) );
  DFFR_X1 \registers_reg[21][25]  ( .D(n3460), .CK(n675), .RN(n6812), .Q(
        \registers[21][25] ) );
  DFFR_X1 \registers_reg[21][24]  ( .D(n3459), .CK(n675), .RN(n6804), .Q(
        \registers[21][24] ) );
  DFFR_X1 \registers_reg[21][23]  ( .D(n3458), .CK(n675), .RN(n6840), .Q(
        \registers[21][23] ) );
  DFFR_X1 \registers_reg[21][22]  ( .D(n3457), .CK(n675), .RN(n6793), .Q(
        \registers[21][22] ) );
  DFFR_X1 \registers_reg[21][21]  ( .D(n3456), .CK(n675), .RN(n6796), .Q(
        \registers[21][21] ) );
  DFFR_X1 \registers_reg[21][20]  ( .D(n3455), .CK(n675), .RN(n6787), .Q(
        \registers[21][20] ) );
  DFFR_X1 \registers_reg[21][19]  ( .D(n3454), .CK(n675), .RN(n6843), .Q(
        \registers[21][19] ) );
  DFFR_X1 \registers_reg[21][18]  ( .D(n3453), .CK(n675), .RN(n6776), .Q(
        \registers[21][18] ) );
  DFFR_X1 \registers_reg[21][17]  ( .D(n3452), .CK(n675), .RN(n6779), .Q(
        \registers[21][17] ) );
  DFFR_X1 \registers_reg[21][16]  ( .D(n3451), .CK(n675), .RN(n6771), .Q(
        \registers[21][16] ) );
  DFFR_X1 \registers_reg[21][15]  ( .D(n3450), .CK(n675), .RN(n6846), .Q(
        \registers[21][15] ) );
  DFFR_X1 \registers_reg[21][14]  ( .D(n3449), .CK(n675), .RN(n6826), .Q(
        \registers[21][14] ) );
  DFFR_X1 \registers_reg[21][13]  ( .D(n3448), .CK(n675), .RN(n6821), .Q(
        \registers[21][13] ) );
  DFFR_X1 \registers_reg[21][12]  ( .D(n3447), .CK(n675), .RN(n6815), .Q(
        \registers[21][12] ) );
  DFFR_X1 \registers_reg[21][11]  ( .D(n3446), .CK(n675), .RN(n6849), .Q(
        \registers[21][11] ) );
  DFFR_X1 \registers_reg[21][10]  ( .D(n3445), .CK(n675), .RN(n6807), .Q(
        \registers[21][10] ) );
  DFFR_X1 \registers_reg[21][9]  ( .D(n3444), .CK(n675), .RN(n6799), .Q(
        \registers[21][9] ) );
  DFFR_X1 \registers_reg[21][8]  ( .D(n3443), .CK(n675), .RN(n6801), .Q(
        \registers[21][8] ) );
  DFFR_X1 \registers_reg[21][7]  ( .D(n3442), .CK(n675), .RN(n6852), .Q(
        \registers[21][7] ) );
  DFFR_X1 \registers_reg[21][6]  ( .D(n3441), .CK(n675), .RN(n6790), .Q(
        \registers[21][6] ) );
  DFFR_X1 \registers_reg[21][5]  ( .D(n3440), .CK(n675), .RN(n6782), .Q(
        \registers[21][5] ) );
  DFFR_X1 \registers_reg[21][4]  ( .D(n3439), .CK(n675), .RN(n6785), .Q(
        \registers[21][4] ) );
  DFFR_X1 \registers_reg[21][3]  ( .D(n3438), .CK(n675), .RN(n6832), .Q(
        \registers[21][3] ) );
  DFFR_X1 \registers_reg[21][2]  ( .D(n3437), .CK(n675), .RN(n6774), .Q(
        \registers[21][2] ) );
  DFFR_X1 \registers_reg[21][1]  ( .D(n3436), .CK(n675), .RN(n6768), .Q(
        \registers[21][1] ) );
  DFFR_X1 \registers_reg[21][0]  ( .D(n3435), .CK(n675), .RN(n6854), .Q(
        \registers[21][0] ) );
  DFFR_X1 \registers_reg[22][31]  ( .D(n3434), .CK(n675), .RN(n6834), .Q(
        \registers[22][31] ) );
  DFFR_X1 \registers_reg[22][30]  ( .D(n3433), .CK(n675), .RN(n6829), .Q(
        \registers[22][30] ) );
  DFFR_X1 \registers_reg[22][29]  ( .D(n3432), .CK(n675), .RN(n6823), .Q(
        \registers[22][29] ) );
  DFFR_X1 \registers_reg[22][28]  ( .D(n3431), .CK(n675), .RN(n6818), .Q(
        \registers[22][28] ) );
  DFFR_X1 \registers_reg[22][27]  ( .D(n3430), .CK(n675), .RN(n6837), .Q(
        \registers[22][27] ) );
  DFFR_X1 \registers_reg[22][26]  ( .D(n3429), .CK(n675), .RN(n6810), .Q(
        \registers[22][26] ) );
  DFFR_X1 \registers_reg[22][25]  ( .D(n3428), .CK(n675), .RN(n6812), .Q(
        \registers[22][25] ) );
  DFFR_X1 \registers_reg[22][24]  ( .D(n3427), .CK(n675), .RN(n6804), .Q(
        \registers[22][24] ) );
  DFFR_X1 \registers_reg[22][23]  ( .D(n3426), .CK(n675), .RN(n6840), .Q(
        \registers[22][23] ) );
  DFFR_X1 \registers_reg[22][22]  ( .D(n3425), .CK(n675), .RN(n6793), .Q(
        \registers[22][22] ) );
  DFFR_X1 \registers_reg[22][21]  ( .D(n3424), .CK(n675), .RN(n6796), .Q(
        \registers[22][21] ) );
  DFFR_X1 \registers_reg[22][20]  ( .D(n3423), .CK(n675), .RN(n6787), .Q(
        \registers[22][20] ) );
  DFFR_X1 \registers_reg[22][19]  ( .D(n3422), .CK(n675), .RN(n6843), .Q(
        \registers[22][19] ) );
  DFFR_X1 \registers_reg[22][18]  ( .D(n3421), .CK(n675), .RN(n6776), .Q(
        \registers[22][18] ) );
  DFFR_X1 \registers_reg[22][17]  ( .D(n3420), .CK(n675), .RN(n6779), .Q(
        \registers[22][17] ) );
  DFFR_X1 \registers_reg[22][16]  ( .D(n3419), .CK(n675), .RN(n6771), .Q(
        \registers[22][16] ) );
  DFFR_X1 \registers_reg[22][15]  ( .D(n3418), .CK(n675), .RN(n6846), .Q(
        \registers[22][15] ) );
  DFFR_X1 \registers_reg[22][14]  ( .D(n3417), .CK(n675), .RN(n6826), .Q(
        \registers[22][14] ) );
  DFFR_X1 \registers_reg[22][13]  ( .D(n3416), .CK(n675), .RN(n6821), .Q(
        \registers[22][13] ) );
  DFFR_X1 \registers_reg[22][12]  ( .D(n3415), .CK(n675), .RN(n6815), .Q(
        \registers[22][12] ) );
  DFFR_X1 \registers_reg[22][11]  ( .D(n3414), .CK(n675), .RN(n6849), .Q(
        \registers[22][11] ) );
  DFFR_X1 \registers_reg[22][10]  ( .D(n3413), .CK(n675), .RN(n6807), .Q(
        \registers[22][10] ) );
  DFFR_X1 \registers_reg[22][9]  ( .D(n3412), .CK(n675), .RN(n6798), .Q(
        \registers[22][9] ) );
  DFFR_X1 \registers_reg[22][8]  ( .D(n3411), .CK(n675), .RN(n6801), .Q(
        \registers[22][8] ) );
  DFFR_X1 \registers_reg[22][7]  ( .D(n3410), .CK(n675), .RN(n6851), .Q(
        \registers[22][7] ) );
  DFFR_X1 \registers_reg[22][6]  ( .D(n3409), .CK(n675), .RN(n6790), .Q(
        \registers[22][6] ) );
  DFFR_X1 \registers_reg[22][5]  ( .D(n3408), .CK(n675), .RN(n6782), .Q(
        \registers[22][5] ) );
  DFFR_X1 \registers_reg[22][4]  ( .D(n3407), .CK(n675), .RN(n6785), .Q(
        \registers[22][4] ) );
  DFFR_X1 \registers_reg[22][3]  ( .D(n3406), .CK(n675), .RN(n6832), .Q(
        \registers[22][3] ) );
  DFFR_X1 \registers_reg[22][2]  ( .D(n3405), .CK(n675), .RN(n6773), .Q(
        \registers[22][2] ) );
  DFFR_X1 \registers_reg[22][1]  ( .D(n3404), .CK(n675), .RN(n6768), .Q(
        \registers[22][1] ) );
  DFFR_X1 \registers_reg[22][0]  ( .D(n3403), .CK(n675), .RN(n6854), .Q(
        \registers[22][0] ) );
  DFFR_X1 \registers_reg[23][31]  ( .D(n3402), .CK(n675), .RN(n6834), .Q(
        \registers[23][31] ) );
  DFFR_X1 \registers_reg[23][30]  ( .D(n3401), .CK(n675), .RN(n6829), .Q(
        \registers[23][30] ) );
  DFFR_X1 \registers_reg[23][29]  ( .D(n3400), .CK(n675), .RN(n6823), .Q(
        \registers[23][29] ) );
  DFFR_X1 \registers_reg[23][28]  ( .D(n3399), .CK(n675), .RN(n6818), .Q(
        \registers[23][28] ) );
  DFFR_X1 \registers_reg[23][27]  ( .D(n3398), .CK(n675), .RN(n6837), .Q(
        \registers[23][27] ) );
  DFFR_X1 \registers_reg[23][26]  ( .D(n3397), .CK(n675), .RN(n6809), .Q(
        \registers[23][26] ) );
  DFFR_X1 \registers_reg[23][25]  ( .D(n3396), .CK(n675), .RN(n6812), .Q(
        \registers[23][25] ) );
  DFFR_X1 \registers_reg[23][24]  ( .D(n3395), .CK(n675), .RN(n6804), .Q(
        \registers[23][24] ) );
  DFFR_X1 \registers_reg[23][23]  ( .D(n3394), .CK(n675), .RN(n6840), .Q(
        \registers[23][23] ) );
  DFFR_X1 \registers_reg[23][22]  ( .D(n3393), .CK(n675), .RN(n6793), .Q(
        \registers[23][22] ) );
  DFFR_X1 \registers_reg[23][21]  ( .D(n3392), .CK(n675), .RN(n6796), .Q(
        \registers[23][21] ) );
  DFFR_X1 \registers_reg[23][20]  ( .D(n3391), .CK(n675), .RN(n6787), .Q(
        \registers[23][20] ) );
  DFFR_X1 \registers_reg[23][19]  ( .D(n3390), .CK(n675), .RN(n6843), .Q(
        \registers[23][19] ) );
  DFFR_X1 \registers_reg[23][18]  ( .D(n3389), .CK(n675), .RN(n6776), .Q(
        \registers[23][18] ) );
  DFFR_X1 \registers_reg[23][17]  ( .D(n3388), .CK(n675), .RN(n6779), .Q(
        \registers[23][17] ) );
  DFFR_X1 \registers_reg[23][16]  ( .D(n3387), .CK(n675), .RN(n6771), .Q(
        \registers[23][16] ) );
  DFFR_X1 \registers_reg[23][15]  ( .D(n3386), .CK(n675), .RN(n6846), .Q(
        \registers[23][15] ) );
  DFFR_X1 \registers_reg[23][14]  ( .D(n3385), .CK(n675), .RN(n6826), .Q(
        \registers[23][14] ) );
  DFFR_X1 \registers_reg[23][13]  ( .D(n3384), .CK(n675), .RN(n6821), .Q(
        \registers[23][13] ) );
  DFFR_X1 \registers_reg[23][12]  ( .D(n3383), .CK(n675), .RN(n6815), .Q(
        \registers[23][12] ) );
  DFFR_X1 \registers_reg[23][11]  ( .D(n3382), .CK(n675), .RN(n6849), .Q(
        \registers[23][11] ) );
  DFFR_X1 \registers_reg[23][10]  ( .D(n3381), .CK(n675), .RN(n6807), .Q(
        \registers[23][10] ) );
  DFFR_X1 \registers_reg[23][9]  ( .D(n3380), .CK(n675), .RN(n6798), .Q(
        \registers[23][9] ) );
  DFFR_X1 \registers_reg[23][8]  ( .D(n3379), .CK(n675), .RN(n6801), .Q(
        \registers[23][8] ) );
  DFFR_X1 \registers_reg[23][7]  ( .D(n3378), .CK(n675), .RN(n6851), .Q(
        \registers[23][7] ) );
  DFFR_X1 \registers_reg[23][6]  ( .D(n3377), .CK(n675), .RN(n6790), .Q(
        \registers[23][6] ) );
  DFFR_X1 \registers_reg[23][5]  ( .D(n3376), .CK(n675), .RN(n6782), .Q(
        \registers[23][5] ) );
  DFFR_X1 \registers_reg[23][4]  ( .D(n3375), .CK(n675), .RN(n6785), .Q(
        \registers[23][4] ) );
  DFFR_X1 \registers_reg[23][3]  ( .D(n3374), .CK(n675), .RN(n6832), .Q(
        \registers[23][3] ) );
  DFFR_X1 \registers_reg[23][2]  ( .D(n3373), .CK(n675), .RN(n6773), .Q(
        \registers[23][2] ) );
  DFFR_X1 \registers_reg[23][1]  ( .D(n3372), .CK(n675), .RN(n6768), .Q(
        \registers[23][1] ) );
  DFFR_X1 \registers_reg[23][0]  ( .D(n3371), .CK(n675), .RN(n6854), .Q(
        \registers[23][0] ) );
  DFFR_X1 \registers_reg[24][31]  ( .D(n3370), .CK(n675), .RN(n6834), .Q(
        \registers[24][31] ), .QN(n5943) );
  DFFR_X1 \registers_reg[24][30]  ( .D(n3369), .CK(n675), .RN(n6829), .Q(
        \registers[24][30] ), .QN(n5942) );
  DFFR_X1 \registers_reg[24][29]  ( .D(n3368), .CK(n675), .RN(n6823), .Q(
        \registers[24][29] ), .QN(n5941) );
  DFFR_X1 \registers_reg[24][28]  ( .D(n3367), .CK(n675), .RN(n6818), .Q(
        \registers[24][28] ), .QN(n5940) );
  DFFR_X1 \registers_reg[24][27]  ( .D(n3366), .CK(n675), .RN(n6837), .Q(
        \registers[24][27] ), .QN(n5981) );
  DFFR_X1 \registers_reg[24][26]  ( .D(n3365), .CK(n675), .RN(n6809), .Q(
        \registers[24][26] ), .QN(n5980) );
  DFFR_X1 \registers_reg[24][25]  ( .D(n3364), .CK(n675), .RN(n6812), .Q(
        \registers[24][25] ), .QN(n5979) );
  DFFR_X1 \registers_reg[24][24]  ( .D(n3363), .CK(n675), .RN(n6804), .Q(
        \registers[24][24] ), .QN(n5978) );
  DFFR_X1 \registers_reg[24][23]  ( .D(n3362), .CK(n675), .RN(n6840), .Q(
        \registers[24][23] ), .QN(n5977) );
  DFFR_X1 \registers_reg[24][22]  ( .D(n3361), .CK(n675), .RN(n6793), .Q(
        \registers[24][22] ), .QN(n5976) );
  DFFR_X1 \registers_reg[24][21]  ( .D(n3360), .CK(n675), .RN(n6796), .Q(
        \registers[24][21] ), .QN(n5939) );
  DFFR_X1 \registers_reg[24][20]  ( .D(n3359), .CK(n675), .RN(n6787), .Q(
        \registers[24][20] ), .QN(n5938) );
  DFFR_X1 \registers_reg[24][19]  ( .D(n3358), .CK(n675), .RN(n6843), .Q(
        \registers[24][19] ), .QN(n5937) );
  DFFR_X1 \registers_reg[24][18]  ( .D(n3357), .CK(n675), .RN(n6776), .Q(
        \registers[24][18] ), .QN(n5936) );
  DFFR_X1 \registers_reg[24][17]  ( .D(n3356), .CK(n675), .RN(n6779), .Q(
        \registers[24][17] ), .QN(n5935) );
  DFFR_X1 \registers_reg[24][16]  ( .D(n3355), .CK(n675), .RN(n6770), .Q(
        \registers[24][16] ), .QN(n5934) );
  DFFR_X1 \registers_reg[24][15]  ( .D(n3354), .CK(n675), .RN(n6846), .Q(
        \registers[24][15] ), .QN(n5933) );
  DFFR_X1 \registers_reg[24][14]  ( .D(n3353), .CK(n675), .RN(n6826), .Q(
        \registers[24][14] ), .QN(n5932) );
  DFFR_X1 \registers_reg[24][13]  ( .D(n3352), .CK(n675), .RN(n6820), .Q(
        \registers[24][13] ), .QN(n5931) );
  DFFR_X1 \registers_reg[24][12]  ( .D(n3351), .CK(n675), .RN(n6815), .Q(
        \registers[24][12] ), .QN(n5930) );
  DFFR_X1 \registers_reg[24][11]  ( .D(n3350), .CK(n675), .RN(n6848), .Q(
        \registers[24][11] ), .QN(n5929) );
  DFFR_X1 \registers_reg[24][10]  ( .D(n3349), .CK(n675), .RN(n6807), .Q(
        \registers[24][10] ), .QN(n5928) );
  DFFR_X1 \registers_reg[24][9]  ( .D(n3348), .CK(n675), .RN(n6798), .Q(
        \registers[24][9] ), .QN(n5927) );
  DFFR_X1 \registers_reg[24][8]  ( .D(n3347), .CK(n675), .RN(n6801), .Q(
        \registers[24][8] ), .QN(n5926) );
  DFFR_X1 \registers_reg[24][7]  ( .D(n3346), .CK(n675), .RN(n6851), .Q(
        \registers[24][7] ), .QN(n5925) );
  DFFR_X1 \registers_reg[24][6]  ( .D(n3345), .CK(n675), .RN(n6790), .Q(
        \registers[24][6] ), .QN(n5924) );
  DFFR_X1 \registers_reg[24][5]  ( .D(n3344), .CK(n675), .RN(n6782), .Q(
        \registers[24][5] ), .QN(n5923) );
  DFFR_X1 \registers_reg[24][4]  ( .D(n3343), .CK(n675), .RN(n6784), .Q(
        \registers[24][4] ), .QN(n5922) );
  DFFR_X1 \registers_reg[24][3]  ( .D(n3342), .CK(n675), .RN(n6832), .Q(
        \registers[24][3] ), .QN(n5921) );
  DFFR_X1 \registers_reg[24][2]  ( .D(n3341), .CK(n675), .RN(n6773), .Q(
        \registers[24][2] ), .QN(n5920) );
  DFFR_X1 \registers_reg[24][1]  ( .D(n3340), .CK(n675), .RN(n6768), .Q(
        \registers[24][1] ), .QN(n5919) );
  DFFR_X1 \registers_reg[24][0]  ( .D(n3339), .CK(n675), .RN(n6854), .Q(
        \registers[24][0] ), .QN(n5918) );
  DFFR_X1 \registers_reg[25][31]  ( .D(n3338), .CK(n675), .RN(n6834), .Q(
        \registers[25][31] ), .QN(n4245) );
  DFFR_X1 \registers_reg[25][30]  ( .D(n3337), .CK(n675), .RN(n6829), .Q(
        \registers[25][30] ), .QN(n4244) );
  DFFR_X1 \registers_reg[25][29]  ( .D(n3336), .CK(n675), .RN(n6823), .Q(
        \registers[25][29] ), .QN(n4243) );
  DFFR_X1 \registers_reg[25][28]  ( .D(n3335), .CK(n675), .RN(n6818), .Q(
        \registers[25][28] ), .QN(n4242) );
  DFFR_X1 \registers_reg[25][27]  ( .D(n3334), .CK(n675), .RN(n6837), .Q(
        \registers[25][27] ), .QN(n4287) );
  DFFR_X1 \registers_reg[25][26]  ( .D(n3333), .CK(n675), .RN(n6809), .Q(
        \registers[25][26] ), .QN(n4284) );
  DFFR_X1 \registers_reg[25][25]  ( .D(n3332), .CK(n675), .RN(n6812), .Q(
        \registers[25][25] ), .QN(n4283) );
  DFFR_X1 \registers_reg[25][24]  ( .D(n3331), .CK(n675), .RN(n6804), .Q(
        \registers[25][24] ), .QN(n4282) );
  DFFR_X1 \registers_reg[25][23]  ( .D(n3330), .CK(n675), .RN(n6840), .Q(
        \registers[25][23] ), .QN(n4281) );
  DFFR_X1 \registers_reg[25][22]  ( .D(n3329), .CK(n675), .RN(n6793), .Q(
        \registers[25][22] ), .QN(n4280) );
  DFFR_X1 \registers_reg[25][21]  ( .D(n3328), .CK(n675), .RN(n6795), .Q(
        \registers[25][21] ), .QN(n4241) );
  DFFR_X1 \registers_reg[25][20]  ( .D(n3327), .CK(n675), .RN(n6787), .Q(
        \registers[25][20] ), .QN(n4240) );
  DFFR_X1 \registers_reg[25][19]  ( .D(n3326), .CK(n675), .RN(n6843), .Q(
        \registers[25][19] ), .QN(n4239) );
  DFFR_X1 \registers_reg[25][18]  ( .D(n3325), .CK(n675), .RN(n6776), .Q(
        \registers[25][18] ), .QN(n4238) );
  DFFR_X1 \registers_reg[25][17]  ( .D(n3324), .CK(n675), .RN(n6779), .Q(
        \registers[25][17] ), .QN(n4237) );
  DFFR_X1 \registers_reg[25][16]  ( .D(n3323), .CK(n675), .RN(n6770), .Q(
        \registers[25][16] ), .QN(n4236) );
  DFFR_X1 \registers_reg[25][15]  ( .D(n3322), .CK(n675), .RN(n6846), .Q(
        \registers[25][15] ), .QN(n4235) );
  DFFR_X1 \registers_reg[25][14]  ( .D(n3321), .CK(n675), .RN(n6826), .Q(
        \registers[25][14] ), .QN(n4234) );
  DFFR_X1 \registers_reg[25][13]  ( .D(n3320), .CK(n675), .RN(n6820), .Q(
        \registers[25][13] ), .QN(n4233) );
  DFFR_X1 \registers_reg[25][12]  ( .D(n3319), .CK(n675), .RN(n6815), .Q(
        \registers[25][12] ), .QN(n4232) );
  DFFR_X1 \registers_reg[25][11]  ( .D(n3318), .CK(n675), .RN(n6848), .Q(
        \registers[25][11] ), .QN(n4231) );
  DFFR_X1 \registers_reg[25][10]  ( .D(n3317), .CK(n675), .RN(n6807), .Q(
        \registers[25][10] ), .QN(n4230) );
  DFFR_X1 \registers_reg[25][9]  ( .D(n3316), .CK(n675), .RN(n6798), .Q(
        \registers[25][9] ), .QN(n4229) );
  DFFR_X1 \registers_reg[25][8]  ( .D(n3315), .CK(n675), .RN(n6801), .Q(
        \registers[25][8] ), .QN(n4228) );
  DFFR_X1 \registers_reg[25][7]  ( .D(n3314), .CK(n675), .RN(n6851), .Q(
        \registers[25][7] ), .QN(n4227) );
  DFFR_X1 \registers_reg[25][6]  ( .D(n3313), .CK(n675), .RN(n6790), .Q(
        \registers[25][6] ), .QN(n4226) );
  DFFR_X1 \registers_reg[25][5]  ( .D(n3312), .CK(n675), .RN(n6782), .Q(
        \registers[25][5] ), .QN(n4225) );
  DFFR_X1 \registers_reg[25][4]  ( .D(n3311), .CK(n675), .RN(n6784), .Q(
        \registers[25][4] ), .QN(n4224) );
  DFFR_X1 \registers_reg[25][3]  ( .D(n3310), .CK(n675), .RN(n6831), .Q(
        \registers[25][3] ), .QN(n4223) );
  DFFR_X1 \registers_reg[25][2]  ( .D(n3309), .CK(n675), .RN(n6773), .Q(
        \registers[25][2] ), .QN(n4222) );
  DFFR_X1 \registers_reg[25][1]  ( .D(n3308), .CK(n675), .RN(n6768), .Q(
        \registers[25][1] ), .QN(n4221) );
  DFFR_X1 \registers_reg[25][0]  ( .D(n3307), .CK(n675), .RN(n6854), .Q(
        \registers[25][0] ), .QN(n4220) );
  DFFR_X1 \registers_reg[26][31]  ( .D(n3306), .CK(n675), .RN(n6834), .Q(
        \registers[26][31] ), .QN(n5896) );
  DFFR_X1 \registers_reg[26][30]  ( .D(n3305), .CK(n675), .RN(n6829), .Q(
        \registers[26][30] ), .QN(n5894) );
  DFFR_X1 \registers_reg[26][29]  ( .D(n3304), .CK(n675), .RN(n6823), .Q(
        \registers[26][29] ), .QN(n5892) );
  DFFR_X1 \registers_reg[26][28]  ( .D(n3303), .CK(n675), .RN(n6818), .Q(
        \registers[26][28] ), .QN(n5890) );
  DFFR_X1 \registers_reg[26][27]  ( .D(n3302), .CK(n675), .RN(n6837), .Q(
        \registers[26][27] ), .QN(n5910) );
  DFFR_X1 \registers_reg[26][26]  ( .D(n3301), .CK(n675), .RN(n6809), .Q(
        \registers[26][26] ), .QN(n5908) );
  DFFR_X1 \registers_reg[26][25]  ( .D(n3300), .CK(n675), .RN(n6812), .Q(
        \registers[26][25] ), .QN(n5906) );
  DFFR_X1 \registers_reg[26][24]  ( .D(n3299), .CK(n675), .RN(n6804), .Q(
        \registers[26][24] ), .QN(n5904) );
  DFFR_X1 \registers_reg[26][23]  ( .D(n3298), .CK(n675), .RN(n6840), .Q(
        \registers[26][23] ), .QN(n5902) );
  DFFR_X1 \registers_reg[26][22]  ( .D(n3297), .CK(n675), .RN(n6793), .Q(
        \registers[26][22] ), .QN(n5900) );
  DFFR_X1 \registers_reg[26][21]  ( .D(n3296), .CK(n675), .RN(n6795), .Q(
        \registers[26][21] ), .QN(n5899) );
  DFFR_X1 \registers_reg[26][20]  ( .D(n3295), .CK(n675), .RN(n6787), .Q(
        \registers[26][20] ), .QN(n5898) );
  DFFR_X1 \registers_reg[26][19]  ( .D(n3294), .CK(n675), .RN(n6843), .Q(
        \registers[26][19] ), .QN(n5880) );
  DFFR_X1 \registers_reg[26][18]  ( .D(n3293), .CK(n675), .RN(n6776), .Q(
        \registers[26][18] ), .QN(n5878) );
  DFFR_X1 \registers_reg[26][17]  ( .D(n3292), .CK(n675), .RN(n6779), .Q(
        \registers[26][17] ), .QN(n5876) );
  DFFR_X1 \registers_reg[26][16]  ( .D(n3291), .CK(n675), .RN(n6770), .Q(
        \registers[26][16] ), .QN(n5874) );
  DFFR_X1 \registers_reg[26][15]  ( .D(n3290), .CK(n675), .RN(n6845), .Q(
        \registers[26][15] ), .QN(n5872) );
  DFFR_X1 \registers_reg[26][14]  ( .D(n3289), .CK(n675), .RN(n6826), .Q(
        \registers[26][14] ), .QN(n5870) );
  DFFR_X1 \registers_reg[26][13]  ( .D(n3288), .CK(n675), .RN(n6820), .Q(
        \registers[26][13] ), .QN(n5868) );
  DFFR_X1 \registers_reg[26][12]  ( .D(n3287), .CK(n675), .RN(n6815), .Q(
        \registers[26][12] ), .QN(n5866) );
  DFFR_X1 \registers_reg[26][11]  ( .D(n3286), .CK(n675), .RN(n6848), .Q(
        \registers[26][11] ), .QN(n5864) );
  DFFR_X1 \registers_reg[26][10]  ( .D(n3285), .CK(n675), .RN(n6806), .Q(
        \registers[26][10] ), .QN(n5862) );
  DFFR_X1 \registers_reg[26][9]  ( .D(n3284), .CK(n675), .RN(n6798), .Q(
        \registers[26][9] ), .QN(n5860) );
  DFFR_X1 \registers_reg[26][8]  ( .D(n3283), .CK(n675), .RN(n6801), .Q(
        \registers[26][8] ), .QN(n5858) );
  DFFR_X1 \registers_reg[26][7]  ( .D(n3282), .CK(n675), .RN(n6851), .Q(
        \registers[26][7] ), .QN(n5856) );
  DFFR_X1 \registers_reg[26][6]  ( .D(n3281), .CK(n675), .RN(n6790), .Q(
        \registers[26][6] ), .QN(n5854) );
  DFFR_X1 \registers_reg[26][5]  ( .D(n3280), .CK(n675), .RN(n6781), .Q(
        \registers[26][5] ), .QN(n5852) );
  DFFR_X1 \registers_reg[26][4]  ( .D(n3279), .CK(n675), .RN(n6784), .Q(
        \registers[26][4] ), .QN(n5850) );
  DFFR_X1 \registers_reg[26][3]  ( .D(n3278), .CK(n675), .RN(n6831), .Q(
        \registers[26][3] ), .QN(n5848) );
  DFFR_X1 \registers_reg[26][2]  ( .D(n3277), .CK(n675), .RN(n6773), .Q(
        \registers[26][2] ), .QN(n5846) );
  DFFR_X1 \registers_reg[26][1]  ( .D(n3276), .CK(n675), .RN(n6768), .Q(
        \registers[26][1] ), .QN(n5844) );
  DFFR_X1 \registers_reg[26][0]  ( .D(n3275), .CK(n675), .RN(n6854), .Q(
        \registers[26][0] ), .QN(n5842) );
  DFFR_X1 \registers_reg[27][31]  ( .D(n3274), .CK(n675), .RN(n6834), .Q(
        \registers[27][31] ), .QN(n4197) );
  DFFR_X1 \registers_reg[27][30]  ( .D(n3273), .CK(n675), .RN(n6828), .Q(
        \registers[27][30] ), .QN(n4195) );
  DFFR_X1 \registers_reg[27][29]  ( .D(n3272), .CK(n675), .RN(n6823), .Q(
        \registers[27][29] ), .QN(n4193) );
  DFFR_X1 \registers_reg[27][28]  ( .D(n3271), .CK(n675), .RN(n6817), .Q(
        \registers[27][28] ), .QN(n4191) );
  DFFR_X1 \registers_reg[27][27]  ( .D(n3270), .CK(n675), .RN(n6837), .Q(
        \registers[27][27] ), .QN(n4211) );
  DFFR_X1 \registers_reg[27][26]  ( .D(n3269), .CK(n675), .RN(n6809), .Q(
        \registers[27][26] ), .QN(n4209) );
  DFFR_X1 \registers_reg[27][25]  ( .D(n3268), .CK(n675), .RN(n6812), .Q(
        \registers[27][25] ), .QN(n4207) );
  DFFR_X1 \registers_reg[27][24]  ( .D(n3267), .CK(n675), .RN(n6804), .Q(
        \registers[27][24] ), .QN(n4205) );
  DFFR_X1 \registers_reg[27][23]  ( .D(n3266), .CK(n675), .RN(n6840), .Q(
        \registers[27][23] ), .QN(n4203) );
  DFFR_X1 \registers_reg[27][22]  ( .D(n3265), .CK(n675), .RN(n6792), .Q(
        \registers[27][22] ), .QN(n4201) );
  DFFR_X1 \registers_reg[27][21]  ( .D(n3264), .CK(n675), .RN(n6795), .Q(
        \registers[27][21] ), .QN(n4200) );
  DFFR_X1 \registers_reg[27][20]  ( .D(n3263), .CK(n675), .RN(n6787), .Q(
        \registers[27][20] ), .QN(n4199) );
  DFFR_X1 \registers_reg[27][19]  ( .D(n3262), .CK(n675), .RN(n6843), .Q(
        \registers[27][19] ), .QN(n4178) );
  DFFR_X1 \registers_reg[27][18]  ( .D(n3261), .CK(n675), .RN(n6776), .Q(
        \registers[27][18] ), .QN(n4176) );
  DFFR_X1 \registers_reg[27][17]  ( .D(n3260), .CK(n675), .RN(n6779), .Q(
        \registers[27][17] ), .QN(n4174) );
  DFFR_X1 \registers_reg[27][16]  ( .D(n3259), .CK(n675), .RN(n6770), .Q(
        \registers[27][16] ), .QN(n4172) );
  DFFR_X1 \registers_reg[27][15]  ( .D(n3258), .CK(n675), .RN(n6845), .Q(
        \registers[27][15] ), .QN(n4170) );
  DFFR_X1 \registers_reg[27][14]  ( .D(n3257), .CK(n675), .RN(n6826), .Q(
        \registers[27][14] ), .QN(n4168) );
  DFFR_X1 \registers_reg[27][13]  ( .D(n3256), .CK(n675), .RN(n6820), .Q(
        \registers[27][13] ), .QN(n4166) );
  DFFR_X1 \registers_reg[27][12]  ( .D(n3255), .CK(n675), .RN(n6815), .Q(
        \registers[27][12] ), .QN(n4164) );
  DFFR_X1 \registers_reg[27][11]  ( .D(n3254), .CK(n675), .RN(n6848), .Q(
        \registers[27][11] ), .QN(n4162) );
  DFFR_X1 \registers_reg[27][10]  ( .D(n3253), .CK(n675), .RN(n6806), .Q(
        \registers[27][10] ), .QN(n4160) );
  DFFR_X1 \registers_reg[27][9]  ( .D(n3252), .CK(n675), .RN(n6798), .Q(
        \registers[27][9] ), .QN(n4158) );
  DFFR_X1 \registers_reg[27][8]  ( .D(n3251), .CK(n675), .RN(n6801), .Q(
        \registers[27][8] ), .QN(n4156) );
  DFFR_X1 \registers_reg[27][7]  ( .D(n3250), .CK(n675), .RN(n6851), .Q(
        \registers[27][7] ), .QN(n4154) );
  DFFR_X1 \registers_reg[27][6]  ( .D(n3249), .CK(n675), .RN(n6790), .Q(
        \registers[27][6] ), .QN(n4152) );
  DFFR_X1 \registers_reg[27][5]  ( .D(n3248), .CK(n675), .RN(n6781), .Q(
        \registers[27][5] ), .QN(n4150) );
  DFFR_X1 \registers_reg[27][4]  ( .D(n3247), .CK(n675), .RN(n6784), .Q(
        \registers[27][4] ), .QN(n2929) );
  DFFR_X1 \registers_reg[27][3]  ( .D(n3246), .CK(n675), .RN(n6831), .Q(
        \registers[27][3] ), .QN(n2860) );
  DFFR_X1 \registers_reg[27][2]  ( .D(n3245), .CK(n675), .RN(n6773), .Q(
        \registers[27][2] ), .QN(n2856) );
  DFFR_X1 \registers_reg[27][1]  ( .D(n3244), .CK(n675), .RN(n6767), .Q(
        \registers[27][1] ), .QN(n2854) );
  DFFR_X1 \registers_reg[27][0]  ( .D(n3243), .CK(n675), .RN(n6854), .Q(
        \registers[27][0] ), .QN(n2852) );
  DFFR_X1 \registers_reg[28][31]  ( .D(n3242), .CK(n675), .RN(n6834), .Q(
        \registers[28][31] ), .QN(n5975) );
  DFFR_X1 \registers_reg[28][30]  ( .D(n3241), .CK(n675), .RN(n6828), .Q(
        \registers[28][30] ), .QN(n5974) );
  DFFR_X1 \registers_reg[28][29]  ( .D(n3240), .CK(n675), .RN(n6823), .Q(
        \registers[28][29] ), .QN(n5973) );
  DFFR_X1 \registers_reg[28][28]  ( .D(n3239), .CK(n675), .RN(n6817), .Q(
        \registers[28][28] ), .QN(n5972) );
  DFFR_X1 \registers_reg[28][27]  ( .D(n3238), .CK(n675), .RN(n6837), .Q(
        \registers[28][27] ), .QN(n5971) );
  DFFR_X1 \registers_reg[28][26]  ( .D(n3237), .CK(n675), .RN(n6809), .Q(
        \registers[28][26] ), .QN(n5970) );
  DFFR_X1 \registers_reg[28][25]  ( .D(n3236), .CK(n675), .RN(n6812), .Q(
        \registers[28][25] ), .QN(n5969) );
  DFFR_X1 \registers_reg[28][24]  ( .D(n3235), .CK(n675), .RN(n6804), .Q(
        \registers[28][24] ), .QN(n5968) );
  DFFR_X1 \registers_reg[28][23]  ( .D(n3234), .CK(n675), .RN(n6840), .Q(
        \registers[28][23] ), .QN(n5967) );
  DFFR_X1 \registers_reg[28][22]  ( .D(n3233), .CK(n675), .RN(n6792), .Q(
        \registers[28][22] ), .QN(n5966) );
  DFFR_X1 \registers_reg[28][21]  ( .D(n3232), .CK(n675), .RN(n6795), .Q(
        \registers[28][21] ), .QN(n5965) );
  DFFR_X1 \registers_reg[28][20]  ( .D(n3231), .CK(n675), .RN(n6787), .Q(
        \registers[28][20] ), .QN(n5964) );
  DFFR_X1 \registers_reg[28][19]  ( .D(n3230), .CK(n675), .RN(n6842), .Q(
        \registers[28][19] ), .QN(n5963) );
  DFFR_X1 \registers_reg[28][18]  ( .D(n3229), .CK(n675), .RN(n6776), .Q(
        \registers[28][18] ), .QN(n5962) );
  DFFR_X1 \registers_reg[28][17]  ( .D(n3228), .CK(n675), .RN(n6779), .Q(
        \registers[28][17] ), .QN(n5961) );
  DFFR_X1 \registers_reg[28][16]  ( .D(n3227), .CK(n675), .RN(n6770), .Q(
        \registers[28][16] ), .QN(n5960) );
  DFFR_X1 \registers_reg[28][15]  ( .D(n3226), .CK(n675), .RN(n6845), .Q(
        \registers[28][15] ), .QN(n5959) );
  DFFR_X1 \registers_reg[28][14]  ( .D(n3225), .CK(n675), .RN(n6826), .Q(
        \registers[28][14] ), .QN(n5958) );
  DFFR_X1 \registers_reg[28][13]  ( .D(n3224), .CK(n675), .RN(n6820), .Q(
        \registers[28][13] ), .QN(n5957) );
  DFFR_X1 \registers_reg[28][12]  ( .D(n3223), .CK(n675), .RN(n6815), .Q(
        \registers[28][12] ), .QN(n5956) );
  DFFR_X1 \registers_reg[28][11]  ( .D(n3222), .CK(n675), .RN(n6848), .Q(
        \registers[28][11] ), .QN(n5955) );
  DFFR_X1 \registers_reg[28][10]  ( .D(n3221), .CK(n675), .RN(n6806), .Q(
        \registers[28][10] ), .QN(n5954) );
  DFFR_X1 \registers_reg[28][9]  ( .D(n3220), .CK(n675), .RN(n6798), .Q(
        \registers[28][9] ), .QN(n5953) );
  DFFR_X1 \registers_reg[28][8]  ( .D(n3219), .CK(n675), .RN(n6801), .Q(
        \registers[28][8] ), .QN(n5952) );
  DFFR_X1 \registers_reg[28][7]  ( .D(n3218), .CK(n675), .RN(n6851), .Q(
        \registers[28][7] ), .QN(n5951) );
  DFFR_X1 \registers_reg[28][6]  ( .D(n3217), .CK(n675), .RN(n6790), .Q(
        \registers[28][6] ), .QN(n5950) );
  DFFR_X1 \registers_reg[28][5]  ( .D(n3216), .CK(n675), .RN(n6781), .Q(
        \registers[28][5] ), .QN(n5949) );
  DFFR_X1 \registers_reg[28][4]  ( .D(n3215), .CK(n675), .RN(n6784), .Q(
        \registers[28][4] ), .QN(n5948) );
  DFFR_X1 \registers_reg[28][3]  ( .D(n3214), .CK(n675), .RN(n6831), .Q(
        \registers[28][3] ), .QN(n5947) );
  DFFR_X1 \registers_reg[28][2]  ( .D(n3213), .CK(n675), .RN(n6773), .Q(
        \registers[28][2] ), .QN(n5946) );
  DFFR_X1 \registers_reg[28][1]  ( .D(n3212), .CK(n675), .RN(n6767), .Q(
        \registers[28][1] ), .QN(n5945) );
  DFFR_X1 \registers_reg[28][0]  ( .D(n3211), .CK(n675), .RN(n6854), .Q(
        \registers[28][0] ), .QN(n5944) );
  DFFR_X1 \registers_reg[29][31]  ( .D(n3210), .CK(n675), .RN(n6834), .Q(
        \registers[29][31] ), .QN(n4279) );
  DFFR_X1 \registers_reg[29][30]  ( .D(n3209), .CK(n675), .RN(n6828), .Q(
        \registers[29][30] ), .QN(n4278) );
  DFFR_X1 \registers_reg[29][29]  ( .D(n3208), .CK(n675), .RN(n6823), .Q(
        \registers[29][29] ), .QN(n4277) );
  DFFR_X1 \registers_reg[29][28]  ( .D(n3207), .CK(n675), .RN(n6817), .Q(
        \registers[29][28] ), .QN(n4276) );
  DFFR_X1 \registers_reg[29][27]  ( .D(n3206), .CK(n675), .RN(n6837), .Q(
        \registers[29][27] ), .QN(n4275) );
  DFFR_X1 \registers_reg[29][26]  ( .D(n3205), .CK(n675), .RN(n6809), .Q(
        \registers[29][26] ), .QN(n4274) );
  DFFR_X1 \registers_reg[29][25]  ( .D(n3204), .CK(n675), .RN(n6812), .Q(
        \registers[29][25] ), .QN(n4273) );
  DFFR_X1 \registers_reg[29][24]  ( .D(n3203), .CK(n675), .RN(n6803), .Q(
        \registers[29][24] ), .QN(n4272) );
  DFFR_X1 \registers_reg[29][23]  ( .D(n3202), .CK(n675), .RN(n6840), .Q(
        \registers[29][23] ), .QN(n4271) );
  DFFR_X1 \registers_reg[29][22]  ( .D(n3201), .CK(n675), .RN(n6792), .Q(
        \registers[29][22] ), .QN(n4270) );
  DFFR_X1 \registers_reg[29][21]  ( .D(n3200), .CK(n675), .RN(n6795), .Q(
        \registers[29][21] ), .QN(n4269) );
  DFFR_X1 \registers_reg[29][20]  ( .D(n3199), .CK(n675), .RN(n6787), .Q(
        \registers[29][20] ), .QN(n4268) );
  DFFR_X1 \registers_reg[29][19]  ( .D(n3198), .CK(n675), .RN(n6842), .Q(
        \registers[29][19] ), .QN(n4267) );
  DFFR_X1 \registers_reg[29][18]  ( .D(n3197), .CK(n675), .RN(n6776), .Q(
        \registers[29][18] ), .QN(n4266) );
  DFFR_X1 \registers_reg[29][17]  ( .D(n3196), .CK(n675), .RN(n6778), .Q(
        \registers[29][17] ), .QN(n4265) );
  DFFR_X1 \registers_reg[29][16]  ( .D(n3195), .CK(n675), .RN(n6770), .Q(
        \registers[29][16] ), .QN(n4264) );
  DFFR_X1 \registers_reg[29][15]  ( .D(n3194), .CK(n675), .RN(n6845), .Q(
        \registers[29][15] ), .QN(n4263) );
  DFFR_X1 \registers_reg[29][14]  ( .D(n3193), .CK(n675), .RN(n6826), .Q(
        \registers[29][14] ), .QN(n4262) );
  DFFR_X1 \registers_reg[29][13]  ( .D(n3192), .CK(n675), .RN(n6820), .Q(
        \registers[29][13] ), .QN(n4261) );
  DFFR_X1 \registers_reg[29][12]  ( .D(n3191), .CK(n675), .RN(n6815), .Q(
        \registers[29][12] ), .QN(n4260) );
  DFFR_X1 \registers_reg[29][11]  ( .D(n3190), .CK(n675), .RN(n6848), .Q(
        \registers[29][11] ), .QN(n4259) );
  DFFR_X1 \registers_reg[29][10]  ( .D(n3189), .CK(n675), .RN(n6806), .Q(
        \registers[29][10] ), .QN(n4258) );
  DFFR_X1 \registers_reg[29][9]  ( .D(n3188), .CK(n675), .RN(n6798), .Q(
        \registers[29][9] ), .QN(n4257) );
  DFFR_X1 \registers_reg[29][8]  ( .D(n3187), .CK(n675), .RN(n6801), .Q(
        \registers[29][8] ), .QN(n4256) );
  DFFR_X1 \registers_reg[29][7]  ( .D(n3186), .CK(n675), .RN(n6851), .Q(
        \registers[29][7] ), .QN(n4255) );
  DFFR_X1 \registers_reg[29][6]  ( .D(n3185), .CK(n675), .RN(n6790), .Q(
        \registers[29][6] ), .QN(n4254) );
  DFFR_X1 \registers_reg[29][5]  ( .D(n3184), .CK(n675), .RN(n6781), .Q(
        \registers[29][5] ), .QN(n4253) );
  DFFR_X1 \registers_reg[29][4]  ( .D(n3183), .CK(n675), .RN(n6784), .Q(
        \registers[29][4] ), .QN(n4250) );
  DFFR_X1 \registers_reg[29][3]  ( .D(n3182), .CK(n675), .RN(n6831), .Q(
        \registers[29][3] ), .QN(n4249) );
  DFFR_X1 \registers_reg[29][2]  ( .D(n3181), .CK(n675), .RN(n6773), .Q(
        \registers[29][2] ), .QN(n4248) );
  DFFR_X1 \registers_reg[29][1]  ( .D(n3180), .CK(n675), .RN(n6767), .Q(
        \registers[29][1] ), .QN(n4247) );
  DFFR_X1 \registers_reg[29][0]  ( .D(n3179), .CK(n675), .RN(n6854), .Q(
        \registers[29][0] ), .QN(n4246) );
  DFFR_X1 \registers_reg[30][31]  ( .D(n3178), .CK(n675), .RN(n6834), .Q(
        \registers[30][31] ) );
  DFFR_X1 \registers_reg[30][30]  ( .D(n3177), .CK(n675), .RN(n6828), .Q(
        \registers[30][30] ) );
  DFFR_X1 \registers_reg[30][29]  ( .D(n3176), .CK(n675), .RN(n6823), .Q(
        \registers[30][29] ) );
  DFFR_X1 \registers_reg[30][28]  ( .D(n3175), .CK(n675), .RN(n6817), .Q(
        \registers[30][28] ) );
  DFFR_X1 \registers_reg[30][27]  ( .D(n3174), .CK(n675), .RN(n6837), .Q(
        \registers[30][27] ) );
  DFFR_X1 \registers_reg[30][26]  ( .D(n3173), .CK(n675), .RN(n6809), .Q(
        \registers[30][26] ) );
  DFFR_X1 \registers_reg[30][25]  ( .D(n3172), .CK(n675), .RN(n6812), .Q(
        \registers[30][25] ) );
  DFFR_X1 \registers_reg[30][24]  ( .D(n3171), .CK(n675), .RN(n6803), .Q(
        \registers[30][24] ) );
  DFFR_X1 \registers_reg[30][23]  ( .D(n3170), .CK(n675), .RN(n6839), .Q(
        \registers[30][23] ) );
  DFFR_X1 \registers_reg[30][22]  ( .D(n3169), .CK(n675), .RN(n6792), .Q(
        \registers[30][22] ) );
  DFFR_X1 \registers_reg[30][21]  ( .D(n3168), .CK(n675), .RN(n6795), .Q(
        \registers[30][21] ) );
  DFFR_X1 \registers_reg[30][20]  ( .D(n3167), .CK(n675), .RN(n6787), .Q(
        \registers[30][20] ) );
  DFFR_X1 \registers_reg[30][19]  ( .D(n3166), .CK(n675), .RN(n6842), .Q(
        \registers[30][19] ) );
  DFFR_X1 \registers_reg[30][18]  ( .D(n3165), .CK(n675), .RN(n6776), .Q(
        \registers[30][18] ) );
  DFFR_X1 \registers_reg[30][17]  ( .D(n3164), .CK(n675), .RN(n6778), .Q(
        \registers[30][17] ) );
  DFFR_X1 \registers_reg[30][16]  ( .D(n3163), .CK(n675), .RN(n6770), .Q(
        \registers[30][16] ) );
  DFFR_X1 \registers_reg[30][15]  ( .D(n3162), .CK(n675), .RN(n6845), .Q(
        \registers[30][15] ) );
  DFFR_X1 \registers_reg[30][14]  ( .D(n3161), .CK(n675), .RN(n6825), .Q(
        \registers[30][14] ) );
  DFFR_X1 \registers_reg[30][13]  ( .D(n3160), .CK(n675), .RN(n6820), .Q(
        \registers[30][13] ) );
  DFFR_X1 \registers_reg[30][12]  ( .D(n3159), .CK(n675), .RN(n6814), .Q(
        \registers[30][12] ) );
  DFFR_X1 \registers_reg[30][11]  ( .D(n3158), .CK(n675), .RN(n6848), .Q(
        \registers[30][11] ) );
  DFFR_X1 \registers_reg[30][10]  ( .D(n3157), .CK(n675), .RN(n6806), .Q(
        \registers[30][10] ) );
  DFFR_X1 \registers_reg[30][9]  ( .D(n3156), .CK(n675), .RN(n6798), .Q(
        \registers[30][9] ) );
  DFFR_X1 \registers_reg[30][8]  ( .D(n3155), .CK(n675), .RN(n6801), .Q(
        \registers[30][8] ) );
  DFFR_X1 \registers_reg[30][7]  ( .D(n3154), .CK(n675), .RN(n6851), .Q(
        \registers[30][7] ) );
  DFFR_X1 \registers_reg[30][6]  ( .D(n3153), .CK(n675), .RN(n6789), .Q(
        \registers[30][6] ) );
  DFFR_X1 \registers_reg[30][5]  ( .D(n3152), .CK(n675), .RN(n6781), .Q(
        \registers[30][5] ) );
  DFFR_X1 \registers_reg[30][4]  ( .D(n3151), .CK(n675), .RN(n6784), .Q(
        \registers[30][4] ) );
  DFFR_X1 \registers_reg[30][3]  ( .D(n3150), .CK(n675), .RN(n6831), .Q(
        \registers[30][3] ) );
  DFFR_X1 \registers_reg[30][2]  ( .D(n3149), .CK(n675), .RN(n6773), .Q(
        \registers[30][2] ) );
  DFFR_X1 \registers_reg[30][1]  ( .D(n3148), .CK(n675), .RN(n6767), .Q(
        \registers[30][1] ) );
  DFFR_X1 \registers_reg[30][0]  ( .D(n3147), .CK(n675), .RN(n6854), .Q(
        \registers[30][0] ) );
  DFFR_X1 \registers_reg[31][31]  ( .D(n3146), .CK(n675), .RN(n6834), .Q(
        \registers[31][31] ) );
  DFFR_X1 \out2_reg[31]  ( .D(n3145), .CK(n675), .RN(n6766), .Q(out2[31]), 
        .QN(n2956) );
  DFFR_X1 \registers_reg[31][30]  ( .D(n3144), .CK(n675), .RN(n6828), .Q(
        \registers[31][30] ) );
  DFFR_X1 \out2_reg[30]  ( .D(n3143), .CK(n675), .RN(n6766), .Q(out2[30]), 
        .QN(n2958) );
  DFFR_X1 \registers_reg[31][29]  ( .D(n3142), .CK(n675), .RN(n6823), .Q(
        \registers[31][29] ) );
  DFFR_X1 \out2_reg[29]  ( .D(n3141), .CK(n675), .RN(n6766), .Q(out2[29]), 
        .QN(n2960) );
  DFFR_X1 \registers_reg[31][28]  ( .D(n3140), .CK(n675), .RN(n6817), .Q(
        \registers[31][28] ) );
  DFFR_X1 \out2_reg[28]  ( .D(n3139), .CK(n675), .RN(n6766), .Q(out2[28]), 
        .QN(n2962) );
  DFFR_X1 \registers_reg[31][27]  ( .D(n3138), .CK(n675), .RN(n6837), .Q(
        \registers[31][27] ) );
  DFFR_X1 \out2_reg[27]  ( .D(n3137), .CK(n675), .RN(n6836), .Q(out2[27]), 
        .QN(n2964) );
  DFFR_X1 \registers_reg[31][26]  ( .D(n3136), .CK(n675), .RN(n6809), .Q(
        \registers[31][26] ) );
  DFFR_X1 \out2_reg[26]  ( .D(n3135), .CK(n675), .RN(n6766), .Q(out2[26]), 
        .QN(n2966) );
  DFFR_X1 \registers_reg[31][25]  ( .D(n3134), .CK(n675), .RN(n6812), .Q(
        \registers[31][25] ) );
  DFFR_X1 \out2_reg[25]  ( .D(n3133), .CK(n675), .RN(n6811), .Q(out2[25]), 
        .QN(n2968) );
  DFFR_X1 \registers_reg[31][24]  ( .D(n3132), .CK(n675), .RN(n6803), .Q(
        \registers[31][24] ) );
  DFFR_X1 \out2_reg[24]  ( .D(n3131), .CK(n675), .RN(n6766), .Q(out2[24]), 
        .QN(n2970) );
  DFFR_X1 \registers_reg[31][23]  ( .D(n3130), .CK(n675), .RN(n6839), .Q(
        \registers[31][23] ) );
  DFFR_X1 \out2_reg[23]  ( .D(n3129), .CK(n675), .RN(n6839), .Q(out2[23]), 
        .QN(n2972) );
  DFFR_X1 \registers_reg[31][22]  ( .D(n3128), .CK(n675), .RN(n6792), .Q(
        \registers[31][22] ) );
  DFFR_X1 \out2_reg[22]  ( .D(n3127), .CK(n675), .RN(n6766), .Q(out2[22]), 
        .QN(n2974) );
  DFFR_X1 \registers_reg[31][21]  ( .D(n3126), .CK(n675), .RN(n6795), .Q(
        \registers[31][21] ) );
  DFFR_X1 \out2_reg[21]  ( .D(n3125), .CK(n675), .RN(n6795), .Q(out2[21]), 
        .QN(n2976) );
  DFFR_X1 \registers_reg[31][20]  ( .D(n3124), .CK(n675), .RN(n6787), .Q(
        \registers[31][20] ) );
  DFFR_X1 \out2_reg[20]  ( .D(n3123), .CK(n675), .RN(n6767), .Q(out2[20]), 
        .QN(n2978) );
  DFFR_X1 \registers_reg[31][19]  ( .D(n3122), .CK(n675), .RN(n6842), .Q(
        \registers[31][19] ) );
  DFFR_X1 \out2_reg[19]  ( .D(n3121), .CK(n675), .RN(n6842), .Q(out2[19]), 
        .QN(n2980) );
  DFFR_X1 \registers_reg[31][18]  ( .D(n3120), .CK(n675), .RN(n6775), .Q(
        \registers[31][18] ) );
  DFFR_X1 \out2_reg[18]  ( .D(n3119), .CK(n675), .RN(n6767), .Q(out2[18]), 
        .QN(n2982) );
  DFFR_X1 \registers_reg[31][17]  ( .D(n3118), .CK(n675), .RN(n6778), .Q(
        \registers[31][17] ) );
  DFFR_X1 \out2_reg[17]  ( .D(n3117), .CK(n675), .RN(n6778), .Q(out2[17]), 
        .QN(n2984) );
  DFFR_X1 \registers_reg[31][16]  ( .D(n3116), .CK(n675), .RN(n6770), .Q(
        \registers[31][16] ) );
  DFFR_X1 \out2_reg[16]  ( .D(n3115), .CK(n675), .RN(n6767), .Q(out2[16]), 
        .QN(n2986) );
  DFFR_X1 \registers_reg[31][15]  ( .D(n3114), .CK(n675), .RN(n6845), .Q(
        \registers[31][15] ) );
  DFFR_X1 \out2_reg[15]  ( .D(n3113), .CK(n675), .RN(n6845), .Q(out2[15]), 
        .QN(n2988) );
  DFFR_X1 \registers_reg[31][14]  ( .D(n3112), .CK(n675), .RN(n6825), .Q(
        \registers[31][14] ) );
  DFFR_X1 \out2_reg[14]  ( .D(n3111), .CK(n675), .RN(n6766), .Q(out2[14]), 
        .QN(n2990) );
  DFFR_X1 \registers_reg[31][13]  ( .D(n3110), .CK(n675), .RN(n6820), .Q(
        \registers[31][13] ) );
  DFFR_X1 \out2_reg[13]  ( .D(n3109), .CK(n675), .RN(n6766), .Q(out2[13]), 
        .QN(n2992) );
  DFFR_X1 \registers_reg[31][12]  ( .D(n3108), .CK(n675), .RN(n6814), .Q(
        \registers[31][12] ) );
  DFFR_X1 \out2_reg[12]  ( .D(n3107), .CK(n675), .RN(n6766), .Q(out2[12]), 
        .QN(n2994) );
  DFFR_X1 \registers_reg[31][11]  ( .D(n3106), .CK(n675), .RN(n6848), .Q(
        \registers[31][11] ) );
  DFFR_X1 \out2_reg[11]  ( .D(n3105), .CK(n675), .RN(n6848), .Q(out2[11]), 
        .QN(n2996) );
  DFFR_X1 \registers_reg[31][10]  ( .D(n3104), .CK(n675), .RN(n6806), .Q(
        \registers[31][10] ) );
  DFFR_X1 \out2_reg[10]  ( .D(n3103), .CK(n675), .RN(n6766), .Q(out2[10]), 
        .QN(n2998) );
  DFFR_X1 \registers_reg[31][9]  ( .D(n3102), .CK(n675), .RN(n6798), .Q(
        \registers[31][9] ) );
  DFFR_X1 \out2_reg[9]  ( .D(n3101), .CK(n675), .RN(n6766), .Q(out2[9]), .QN(
        n3000) );
  DFFR_X1 \registers_reg[31][8]  ( .D(n3100), .CK(n675), .RN(n6801), .Q(
        \registers[31][8] ) );
  DFFR_X1 \out2_reg[8]  ( .D(n3099), .CK(n675), .RN(n6800), .Q(out2[8]), .QN(
        n3002) );
  DFFR_X1 \registers_reg[31][7]  ( .D(n3098), .CK(n675), .RN(n6851), .Q(
        \registers[31][7] ) );
  DFFR_X1 \out2_reg[7]  ( .D(n3097), .CK(n675), .RN(n6851), .Q(out2[7]), .QN(
        n3004) );
  DFFR_X1 \registers_reg[31][6]  ( .D(n3096), .CK(n675), .RN(n6789), .Q(
        \registers[31][6] ) );
  DFFR_X1 \out2_reg[6]  ( .D(n3095), .CK(n675), .RN(n6767), .Q(out2[6]), .QN(
        n3006) );
  DFFR_X1 \registers_reg[31][5]  ( .D(n3094), .CK(n675), .RN(n6781), .Q(
        \registers[31][5] ) );
  DFFR_X1 \out2_reg[5]  ( .D(n3093), .CK(n675), .RN(n6767), .Q(out2[5]), .QN(
        n3008) );
  DFFR_X1 \registers_reg[31][4]  ( .D(n3092), .CK(n675), .RN(n6784), .Q(
        \registers[31][4] ) );
  DFFR_X1 \out2_reg[4]  ( .D(n3091), .CK(n675), .RN(n6784), .Q(out2[4]), .QN(
        n3010) );
  DFFR_X1 \registers_reg[31][3]  ( .D(n3090), .CK(n675), .RN(n6831), .Q(
        \registers[31][3] ) );
  DFFR_X1 \out2_reg[3]  ( .D(n3089), .CK(n675), .RN(n6831), .Q(out2[3]), .QN(
        n3012) );
  DFFR_X1 \registers_reg[31][2]  ( .D(n3088), .CK(n675), .RN(n6773), .Q(
        \registers[31][2] ) );
  DFFR_X1 \out2_reg[2]  ( .D(n3087), .CK(n675), .RN(n6773), .Q(out2[2]), .QN(
        n3014) );
  DFFR_X1 \registers_reg[31][1]  ( .D(n3086), .CK(n675), .RN(n6767), .Q(
        \registers[31][1] ) );
  DFFR_X1 \out2_reg[1]  ( .D(n3085), .CK(n675), .RN(n6767), .Q(out2[1]), .QN(
        n3016) );
  DFFR_X1 \registers_reg[31][0]  ( .D(n3084), .CK(n675), .RN(n6854), .Q(
        \registers[31][0] ) );
  DFFR_X1 \out2_reg[0]  ( .D(n3083), .CK(n675), .RN(n6853), .Q(out2[0]), .QN(
        n3018) );
  DFFR_X1 \out1_reg[31]  ( .D(n3082), .CK(n675), .RN(n6834), .Q(out1[31]), 
        .QN(n3019) );
  DFFR_X1 \out1_reg[30]  ( .D(n3081), .CK(n675), .RN(n6828), .Q(out1[30]), 
        .QN(n3020) );
  DFFR_X1 \out1_reg[29]  ( .D(n3080), .CK(n675), .RN(n6823), .Q(out1[29]), 
        .QN(n3021) );
  DFFR_X1 \out1_reg[28]  ( .D(n3079), .CK(n675), .RN(n6817), .Q(out1[28]), 
        .QN(n3022) );
  DFFR_X1 \out1_reg[27]  ( .D(n3078), .CK(n675), .RN(n6836), .Q(out1[27]), 
        .QN(n3023) );
  DFFR_X1 \out1_reg[26]  ( .D(n3077), .CK(n675), .RN(n6809), .Q(out1[26]), 
        .QN(n3024) );
  DFFR_X1 \out1_reg[25]  ( .D(n3076), .CK(n675), .RN(n6812), .Q(out1[25]), 
        .QN(n3025) );
  DFFR_X1 \out1_reg[24]  ( .D(n3075), .CK(n675), .RN(n6803), .Q(out1[24]), 
        .QN(n3026) );
  DFFR_X1 \out1_reg[23]  ( .D(n3074), .CK(n675), .RN(n6839), .Q(out1[23]), 
        .QN(n3027) );
  DFFR_X1 \out1_reg[22]  ( .D(n3073), .CK(n675), .RN(n6792), .Q(out1[22]), 
        .QN(n3028) );
  DFFR_X1 \out1_reg[21]  ( .D(n3072), .CK(n675), .RN(n6795), .Q(out1[21]), 
        .QN(n3029) );
  DFFR_X1 \out1_reg[20]  ( .D(n3071), .CK(n675), .RN(n6787), .Q(out1[20]), 
        .QN(n3030) );
  DFFR_X1 \out1_reg[19]  ( .D(n3070), .CK(n675), .RN(n6842), .Q(out1[19]), 
        .QN(n3031) );
  DFFR_X1 \out1_reg[18]  ( .D(n3069), .CK(n675), .RN(n6775), .Q(out1[18]), 
        .QN(n3032) );
  DFFR_X1 \out1_reg[17]  ( .D(n3068), .CK(n675), .RN(n6778), .Q(out1[17]), 
        .QN(n3033) );
  DFFR_X1 \out1_reg[16]  ( .D(n3067), .CK(n675), .RN(n6770), .Q(out1[16]), 
        .QN(n3034) );
  DFFR_X1 \out1_reg[15]  ( .D(n3066), .CK(n675), .RN(n6845), .Q(out1[15]), 
        .QN(n3035) );
  DFFR_X1 \out1_reg[14]  ( .D(n3065), .CK(n675), .RN(n6825), .Q(out1[14]), 
        .QN(n3036) );
  DFFR_X1 \out1_reg[13]  ( .D(n3064), .CK(n675), .RN(n6820), .Q(out1[13]), 
        .QN(n3037) );
  DFFR_X1 \out1_reg[12]  ( .D(n3063), .CK(n675), .RN(n6814), .Q(out1[12]), 
        .QN(n3038) );
  DFFR_X1 \out1_reg[11]  ( .D(n3062), .CK(n675), .RN(n6848), .Q(out1[11]), 
        .QN(n3039) );
  DFFR_X1 \out1_reg[10]  ( .D(n3061), .CK(n675), .RN(n6806), .Q(out1[10]), 
        .QN(n3040) );
  DFFR_X1 \out1_reg[9]  ( .D(n3060), .CK(n675), .RN(n6798), .Q(out1[9]), .QN(
        n3041) );
  DFFR_X1 \out1_reg[8]  ( .D(n3059), .CK(n675), .RN(n6800), .Q(out1[8]), .QN(
        n3042) );
  DFFR_X1 \out1_reg[7]  ( .D(n3058), .CK(n675), .RN(n6851), .Q(out1[7]), .QN(
        n3043) );
  DFFR_X1 \out1_reg[6]  ( .D(n3057), .CK(n675), .RN(n6789), .Q(out1[6]), .QN(
        n3044) );
  DFFR_X1 \out1_reg[5]  ( .D(n3056), .CK(n675), .RN(n6781), .Q(out1[5]), .QN(
        n3045) );
  DFFR_X1 \out1_reg[4]  ( .D(n3055), .CK(n675), .RN(n6784), .Q(out1[4]), .QN(
        n3046) );
  DFFR_X1 \out1_reg[3]  ( .D(n3054), .CK(n675), .RN(n6831), .Q(out1[3]), .QN(
        n3047) );
  DFFR_X1 \out1_reg[2]  ( .D(n3053), .CK(n675), .RN(n6773), .Q(out1[2]), .QN(
        n3048) );
  DFFR_X1 \out1_reg[1]  ( .D(n3052), .CK(n675), .RN(n6767), .Q(out1[1]), .QN(
        n3049) );
  DFFR_X1 \out1_reg[0]  ( .D(n3051), .CK(n675), .RN(n6853), .Q(out1[0]), .QN(
        n3050) );
  INV_X2 U3 ( .A(clk), .ZN(n675) );
  NOR2_X1 U4 ( .A1(n5751), .A2(add_rd1[2]), .ZN(n5736) );
  NOR3_X1 U5 ( .A1(add_rd1[0]), .A2(add_rd1[4]), .A3(n5744), .ZN(n5729) );
  NOR2_X1 U6 ( .A1(add_rd1[1]), .A2(add_rd1[2]), .ZN(n5724) );
  NOR3_X1 U7 ( .A1(add_rd1[3]), .A2(add_rd1[4]), .A3(n5745), .ZN(n5726) );
  NOR3_X1 U8 ( .A1(add_rd1[3]), .A2(add_rd1[4]), .A3(add_rd1[0]), .ZN(n5725)
         );
  NOR2_X1 U9 ( .A1(n5083), .A2(add_rd2[2]), .ZN(n5068) );
  NOR3_X1 U10 ( .A1(add_rd2[0]), .A2(add_rd2[4]), .A3(n5076), .ZN(n5061) );
  NOR3_X1 U11 ( .A1(n5081), .A2(add_rd2[0]), .A3(n5076), .ZN(n5067) );
  NOR2_X1 U12 ( .A1(n5080), .A2(add_rd2[1]), .ZN(n5059) );
  NOR2_X1 U13 ( .A1(add_rd2[1]), .A2(add_rd2[2]), .ZN(n5056) );
  NOR3_X1 U14 ( .A1(add_rd2[0]), .A2(add_rd2[3]), .A3(n5081), .ZN(n5064) );
  NOR2_X1 U15 ( .A1(n4354), .A2(add_wr[1]), .ZN(n1786) );
  NOR2_X1 U16 ( .A1(add_wr[0]), .A2(add_wr[1]), .ZN(n1750) );
  AND2_X1 U17 ( .A1(n1786), .A2(n1751), .ZN(n2560) );
  BUF_X1 U18 ( .A(n6492), .Z(n5982) );
  BUF_X1 U19 ( .A(n6492), .Z(n5983) );
  BUF_X1 U20 ( .A(n6501), .Z(n5985) );
  BUF_X1 U21 ( .A(n6501), .Z(n5986) );
  BUF_X1 U22 ( .A(n6559), .Z(n6006) );
  BUF_X1 U23 ( .A(n6559), .Z(n6007) );
  BUF_X1 U24 ( .A(n6568), .Z(n6009) );
  BUF_X1 U25 ( .A(n6568), .Z(n6010) );
  BUF_X1 U26 ( .A(n6577), .Z(n6012) );
  BUF_X1 U27 ( .A(n6577), .Z(n6013) );
  BUF_X1 U28 ( .A(n6586), .Z(n6015) );
  BUF_X1 U29 ( .A(n6586), .Z(n6016) );
  BUF_X1 U30 ( .A(n6628), .Z(n6030) );
  BUF_X1 U31 ( .A(n6628), .Z(n6031) );
  BUF_X1 U32 ( .A(n6637), .Z(n6033) );
  BUF_X1 U33 ( .A(n6637), .Z(n6034) );
  BUF_X1 U34 ( .A(n6646), .Z(n6036) );
  BUF_X1 U35 ( .A(n6646), .Z(n6037) );
  BUF_X1 U36 ( .A(n6655), .Z(n6039) );
  BUF_X1 U37 ( .A(n6655), .Z(n6040) );
  BUF_X1 U38 ( .A(n6714), .Z(n6060) );
  BUF_X1 U39 ( .A(n6714), .Z(n6061) );
  BUF_X1 U40 ( .A(n6723), .Z(n6063) );
  BUF_X1 U41 ( .A(n6723), .Z(n6064) );
  BUF_X1 U42 ( .A(n4321), .Z(n5988) );
  BUF_X1 U43 ( .A(n4321), .Z(n5989) );
  BUF_X1 U44 ( .A(n4286), .Z(n5991) );
  BUF_X1 U45 ( .A(n4286), .Z(n5992) );
  BUF_X1 U46 ( .A(n4252), .Z(n5994) );
  BUF_X1 U47 ( .A(n4252), .Z(n5995) );
  BUF_X1 U48 ( .A(n6533), .Z(n5997) );
  BUF_X1 U49 ( .A(n6533), .Z(n5998) );
  BUF_X1 U50 ( .A(n4184), .Z(n6000) );
  BUF_X1 U51 ( .A(n4184), .Z(n6001) );
  BUF_X1 U52 ( .A(n4149), .Z(n6003) );
  BUF_X1 U53 ( .A(n4149), .Z(n6004) );
  BUF_X1 U54 ( .A(n2825), .Z(n6018) );
  BUF_X1 U55 ( .A(n2825), .Z(n6019) );
  BUF_X1 U56 ( .A(n6602), .Z(n6021) );
  BUF_X1 U57 ( .A(n6602), .Z(n6022) );
  BUF_X1 U58 ( .A(n2757), .Z(n6024) );
  BUF_X1 U59 ( .A(n2757), .Z(n6025) );
  BUF_X1 U60 ( .A(n2722), .Z(n6027) );
  BUF_X1 U61 ( .A(n2722), .Z(n6028) );
  BUF_X1 U62 ( .A(n6664), .Z(n6042) );
  BUF_X1 U63 ( .A(n6664), .Z(n6043) );
  BUF_X1 U64 ( .A(n6672), .Z(n6045) );
  BUF_X1 U65 ( .A(n6672), .Z(n6046) );
  BUF_X1 U66 ( .A(n6682), .Z(n6048) );
  BUF_X1 U67 ( .A(n6682), .Z(n6049) );
  BUF_X1 U68 ( .A(n6690), .Z(n6051) );
  BUF_X1 U69 ( .A(n6690), .Z(n6052) );
  BUF_X1 U70 ( .A(n6491), .Z(n5984) );
  BUF_X1 U71 ( .A(n6500), .Z(n5987) );
  BUF_X1 U72 ( .A(n6558), .Z(n6008) );
  BUF_X1 U73 ( .A(n6567), .Z(n6011) );
  BUF_X1 U74 ( .A(n6576), .Z(n6014) );
  BUF_X1 U75 ( .A(n6585), .Z(n6017) );
  BUF_X1 U76 ( .A(n6627), .Z(n6032) );
  BUF_X1 U77 ( .A(n6636), .Z(n6035) );
  BUF_X1 U78 ( .A(n6645), .Z(n6038) );
  BUF_X1 U79 ( .A(n6654), .Z(n6041) );
  BUF_X1 U80 ( .A(n6713), .Z(n6062) );
  BUF_X1 U81 ( .A(n6722), .Z(n6065) );
  BUF_X1 U82 ( .A(n4321), .Z(n5990) );
  BUF_X1 U83 ( .A(n4286), .Z(n5993) );
  BUF_X1 U84 ( .A(n4252), .Z(n5996) );
  BUF_X1 U85 ( .A(n6533), .Z(n5999) );
  BUF_X1 U86 ( .A(n4184), .Z(n6002) );
  BUF_X1 U87 ( .A(n4149), .Z(n6005) );
  BUF_X1 U88 ( .A(n2825), .Z(n6020) );
  BUF_X1 U89 ( .A(n6602), .Z(n6023) );
  BUF_X1 U90 ( .A(n2757), .Z(n6026) );
  BUF_X1 U91 ( .A(n2722), .Z(n6029) );
  BUF_X1 U92 ( .A(n6663), .Z(n6044) );
  BUF_X1 U93 ( .A(n6673), .Z(n6047) );
  BUF_X1 U94 ( .A(n6681), .Z(n6050) );
  BUF_X1 U95 ( .A(n6691), .Z(n6053) );
  AND2_X1 U96 ( .A1(n5069), .A2(n5070), .ZN(n6392) );
  AND2_X1 U97 ( .A1(n5069), .A2(n5070), .ZN(n6391) );
  AND2_X1 U98 ( .A1(n5069), .A2(n5070), .ZN(n4417) );
  BUF_X1 U99 ( .A(n1964), .Z(n6054) );
  BUF_X1 U100 ( .A(n1964), .Z(n6055) );
  BUF_X1 U101 ( .A(n1930), .Z(n6057) );
  BUF_X1 U102 ( .A(n1930), .Z(n6058) );
  INV_X1 U103 ( .A(n6745), .ZN(n6735) );
  INV_X1 U104 ( .A(n6745), .ZN(n6736) );
  BUF_X1 U105 ( .A(n1964), .Z(n6056) );
  BUF_X1 U106 ( .A(n1930), .Z(n6059) );
  BUF_X1 U107 ( .A(n4413), .Z(n6419) );
  BUF_X1 U108 ( .A(n4442), .Z(n6289) );
  BUF_X1 U109 ( .A(n4413), .Z(n6420) );
  BUF_X1 U110 ( .A(n4442), .Z(n6290) );
  BUF_X1 U111 ( .A(n4427), .Z(n6379) );
  BUF_X1 U112 ( .A(n4427), .Z(n6380) );
  BUF_X1 U113 ( .A(n4413), .Z(n6421) );
  BUF_X1 U114 ( .A(n4442), .Z(n6291) );
  BUF_X1 U115 ( .A(n4427), .Z(n6381) );
  INV_X1 U116 ( .A(n4406), .ZN(n6480) );
  INV_X1 U117 ( .A(n4411), .ZN(n6455) );
  INV_X1 U118 ( .A(n4410), .ZN(n6447) );
  INV_X1 U119 ( .A(n4405), .ZN(n6472) );
  INV_X1 U120 ( .A(n4421), .ZN(n6403) );
  INV_X1 U121 ( .A(n4445), .ZN(n6300) );
  INV_X1 U122 ( .A(n4434), .ZN(n6355) );
  INV_X1 U123 ( .A(n4439), .ZN(n6324) );
  INV_X1 U124 ( .A(n4420), .ZN(n6395) );
  INV_X1 U125 ( .A(n4444), .ZN(n6292) );
  INV_X1 U126 ( .A(n4435), .ZN(n6363) );
  BUF_X1 U127 ( .A(n6382), .Z(n6383) );
  BUF_X1 U128 ( .A(n6382), .Z(n6384) );
  BUF_X1 U129 ( .A(n6422), .Z(n6423) );
  BUF_X1 U130 ( .A(n6422), .Z(n6424) );
  BUF_X1 U131 ( .A(n6332), .Z(n6333) );
  BUF_X1 U132 ( .A(n6332), .Z(n6334) );
  BUF_X1 U133 ( .A(n6463), .Z(n6464) );
  BUF_X1 U134 ( .A(n6463), .Z(n6465) );
  BUF_X1 U135 ( .A(n6382), .Z(n6385) );
  BUF_X1 U136 ( .A(n4429), .Z(n6386) );
  BUF_X1 U137 ( .A(n4429), .Z(n6387) );
  BUF_X1 U138 ( .A(n4429), .Z(n6388) );
  BUF_X1 U139 ( .A(n6422), .Z(n6425) );
  BUF_X1 U140 ( .A(n4415), .Z(n6426) );
  BUF_X1 U141 ( .A(n4415), .Z(n6427) );
  BUF_X1 U142 ( .A(n4415), .Z(n6428) );
  BUF_X1 U143 ( .A(n6332), .Z(n6335) );
  BUF_X1 U144 ( .A(n4440), .Z(n6336) );
  BUF_X1 U145 ( .A(n4440), .Z(n6337) );
  BUF_X1 U146 ( .A(n4440), .Z(n6338) );
  BUF_X1 U147 ( .A(n6463), .Z(n6466) );
  BUF_X1 U148 ( .A(n4402), .Z(n6467) );
  BUF_X1 U149 ( .A(n4402), .Z(n6468) );
  BUF_X1 U150 ( .A(n4402), .Z(n6469) );
  INV_X1 U151 ( .A(n6512), .ZN(n4321) );
  INV_X1 U152 ( .A(n6519), .ZN(n4286) );
  INV_X1 U153 ( .A(n6545), .ZN(n4184) );
  INV_X1 U154 ( .A(n6552), .ZN(n4149) );
  INV_X1 U155 ( .A(n6614), .ZN(n2757) );
  INV_X1 U156 ( .A(n6621), .ZN(n2722) );
  INV_X1 U157 ( .A(n6528), .ZN(n4252) );
  INV_X1 U158 ( .A(n6597), .ZN(n2825) );
  BUF_X1 U159 ( .A(n6762), .Z(n6872) );
  BUF_X1 U160 ( .A(n6755), .Z(n6857) );
  BUF_X1 U161 ( .A(n6762), .Z(n6871) );
  BUF_X1 U162 ( .A(n6761), .Z(n6869) );
  BUF_X1 U163 ( .A(n6761), .Z(n6870) );
  BUF_X1 U164 ( .A(n6755), .Z(n6858) );
  BUF_X1 U165 ( .A(n6760), .Z(n6868) );
  BUF_X1 U166 ( .A(n6759), .Z(n6866) );
  BUF_X1 U167 ( .A(n6760), .Z(n6867) );
  BUF_X1 U168 ( .A(n6759), .Z(n6865) );
  BUF_X1 U169 ( .A(n6758), .Z(n6864) );
  BUF_X1 U170 ( .A(n6756), .Z(n6859) );
  BUF_X1 U171 ( .A(n6758), .Z(n6863) );
  BUF_X1 U172 ( .A(n6757), .Z(n6862) );
  BUF_X1 U173 ( .A(n6757), .Z(n6861) );
  BUF_X1 U174 ( .A(n6756), .Z(n6860) );
  NOR3_X1 U175 ( .A1(n5076), .A2(n5081), .A3(n5077), .ZN(n5069) );
  NOR2_X1 U176 ( .A1(n5083), .A2(n5080), .ZN(n5070) );
  NAND2_X1 U177 ( .A1(n5068), .A2(n5061), .ZN(n6389) );
  NAND2_X1 U178 ( .A1(n5068), .A2(n5061), .ZN(n6390) );
  NAND2_X1 U179 ( .A1(n5064), .A2(n5056), .ZN(n6429) );
  NAND2_X1 U180 ( .A1(n5064), .A2(n5056), .ZN(n6430) );
  INV_X1 U181 ( .A(n6754), .ZN(n6746) );
  INV_X1 U182 ( .A(n6754), .ZN(n6747) );
  NAND2_X1 U183 ( .A1(n5068), .A2(n5061), .ZN(n4430) );
  NAND2_X1 U184 ( .A1(n5064), .A2(n5056), .ZN(n4416) );
  AND2_X1 U185 ( .A1(n5067), .A2(n5070), .ZN(n6393) );
  AND2_X1 U186 ( .A1(n5067), .A2(n5070), .ZN(n6394) );
  AND2_X1 U187 ( .A1(n5059), .A2(n5057), .ZN(n6470) );
  AND2_X1 U188 ( .A1(n5059), .A2(n5057), .ZN(n6471) );
  AND2_X1 U189 ( .A1(n5067), .A2(n5070), .ZN(n4418) );
  AND2_X1 U190 ( .A1(n5059), .A2(n5057), .ZN(n4403) );
  BUF_X1 U191 ( .A(n1823), .Z(n6066) );
  BUF_X1 U192 ( .A(n1823), .Z(n6067) );
  BUF_X1 U193 ( .A(n1788), .Z(n6069) );
  BUF_X1 U194 ( .A(n1788), .Z(n6070) );
  NAND2_X1 U195 ( .A1(n5056), .A2(n5061), .ZN(n4411) );
  NAND2_X1 U196 ( .A1(n5056), .A2(n5062), .ZN(n4410) );
  NAND2_X1 U197 ( .A1(n5056), .A2(n5058), .ZN(n4405) );
  NAND2_X1 U198 ( .A1(n5056), .A2(n5057), .ZN(n4406) );
  NAND2_X1 U199 ( .A1(n5067), .A2(n5068), .ZN(n4421) );
  NAND2_X1 U200 ( .A1(n5064), .A2(n5068), .ZN(n4445) );
  NAND2_X1 U201 ( .A1(n5057), .A2(n5068), .ZN(n4434) );
  NAND2_X1 U202 ( .A1(n5069), .A2(n5068), .ZN(n4420) );
  NAND2_X1 U203 ( .A1(n5069), .A2(n5059), .ZN(n4439) );
  NAND2_X1 U204 ( .A1(n5067), .A2(n5059), .ZN(n6332) );
  NAND2_X1 U205 ( .A1(n5067), .A2(n5059), .ZN(n4440) );
  NAND2_X1 U206 ( .A1(n5065), .A2(n5068), .ZN(n4444) );
  NAND2_X1 U207 ( .A1(n5058), .A2(n5068), .ZN(n4435) );
  BUF_X1 U208 ( .A(n1823), .Z(n6068) );
  BUF_X1 U209 ( .A(n1788), .Z(n6071) );
  NAND2_X1 U210 ( .A1(n5062), .A2(n5068), .ZN(n6382) );
  NAND2_X1 U211 ( .A1(n5062), .A2(n5068), .ZN(n4429) );
  NAND2_X1 U212 ( .A1(n5065), .A2(n5056), .ZN(n6422) );
  NAND2_X1 U213 ( .A1(n5065), .A2(n5056), .ZN(n4415) );
  AND2_X1 U214 ( .A1(n5056), .A2(n5067), .ZN(n4437) );
  AND2_X1 U215 ( .A1(n5056), .A2(n5069), .ZN(n4436) );
  AND2_X1 U216 ( .A1(n5059), .A2(n5061), .ZN(n4408) );
  AND2_X1 U217 ( .A1(n5059), .A2(n5062), .ZN(n4407) );
  AND2_X1 U218 ( .A1(n5057), .A2(n5070), .ZN(n4431) );
  AND2_X1 U219 ( .A1(n5070), .A2(n5062), .ZN(n4426) );
  AND2_X1 U220 ( .A1(n5065), .A2(n5059), .ZN(n4412) );
  AND2_X1 U221 ( .A1(n5065), .A2(n5070), .ZN(n4441) );
  AND2_X1 U222 ( .A1(n5058), .A2(n5070), .ZN(n4432) );
  AND2_X1 U223 ( .A1(n5064), .A2(n5059), .ZN(n4413) );
  AND2_X1 U224 ( .A1(n5064), .A2(n5070), .ZN(n4442) );
  AND2_X1 U225 ( .A1(n5059), .A2(n5058), .ZN(n6463) );
  AND2_X1 U226 ( .A1(n5059), .A2(n5058), .ZN(n4402) );
  AND2_X1 U227 ( .A1(n5070), .A2(n5061), .ZN(n4427) );
  BUF_X1 U228 ( .A(n2560), .Z(n6745) );
  BUF_X1 U229 ( .A(n6741), .Z(n6744) );
  BUF_X1 U230 ( .A(n6742), .Z(n6743) );
  BUF_X1 U231 ( .A(n2560), .Z(n6742) );
  BUF_X1 U232 ( .A(n2560), .Z(n6741) );
  BUF_X1 U233 ( .A(n2560), .Z(n6740) );
  BUF_X1 U234 ( .A(n2560), .Z(n6739) );
  BUF_X1 U235 ( .A(n2560), .Z(n6738) );
  BUF_X1 U236 ( .A(n2560), .Z(n6737) );
  INV_X1 U237 ( .A(n6700), .ZN(n1964) );
  INV_X1 U238 ( .A(n6707), .ZN(n1930) );
  BUF_X1 U239 ( .A(n6763), .Z(n6762) );
  BUF_X1 U240 ( .A(n6763), .Z(n6761) );
  BUF_X1 U241 ( .A(n6763), .Z(n6760) );
  BUF_X1 U242 ( .A(n6764), .Z(n6759) );
  BUF_X1 U243 ( .A(n6764), .Z(n6758) );
  BUF_X1 U244 ( .A(n6764), .Z(n6757) );
  BUF_X1 U245 ( .A(n6765), .Z(n6755) );
  BUF_X1 U246 ( .A(n6765), .Z(n6756) );
  NOR3_X1 U247 ( .A1(add_rd2[3]), .A2(add_rd2[4]), .A3(add_rd2[0]), .ZN(n5057)
         );
  NOR3_X1 U248 ( .A1(n5076), .A2(add_rd2[4]), .A3(n5077), .ZN(n5062) );
  NOR3_X1 U249 ( .A1(n5081), .A2(add_rd2[3]), .A3(n5077), .ZN(n5065) );
  NOR3_X1 U250 ( .A1(add_rd2[3]), .A2(add_rd2[4]), .A3(n5077), .ZN(n5058) );
  AND2_X1 U251 ( .A1(n5737), .A2(n5738), .ZN(n6182) );
  AND2_X1 U252 ( .A1(n5737), .A2(n5738), .ZN(n6183) );
  AND2_X1 U253 ( .A1(n5737), .A2(n5738), .ZN(n5116) );
  INV_X1 U254 ( .A(add_rd2[4]), .ZN(n5081) );
  BUF_X1 U255 ( .A(n5131), .Z(n6143) );
  BUF_X1 U256 ( .A(n5131), .Z(n6144) );
  BUF_X1 U257 ( .A(n5107), .Z(n6242) );
  BUF_X1 U258 ( .A(n5136), .Z(n6116) );
  BUF_X1 U259 ( .A(n5126), .Z(n6170) );
  BUF_X1 U260 ( .A(n5107), .Z(n6243) );
  BUF_X1 U261 ( .A(n5136), .Z(n6117) );
  BUF_X1 U262 ( .A(n5126), .Z(n6171) );
  BUF_X1 U263 ( .A(n5131), .Z(n6145) );
  BUF_X1 U264 ( .A(n5107), .Z(n6244) );
  BUF_X1 U265 ( .A(n5136), .Z(n6118) );
  BUF_X1 U266 ( .A(n5126), .Z(n6172) );
  INV_X1 U267 ( .A(add_rd2[0]), .ZN(n5077) );
  INV_X1 U268 ( .A(add_rd2[3]), .ZN(n5076) );
  INV_X1 U269 ( .A(n5133), .ZN(n6146) );
  INV_X1 U270 ( .A(n5110), .ZN(n6253) );
  INV_X1 U271 ( .A(n5109), .ZN(n6245) );
  INV_X1 U272 ( .A(n5134), .ZN(n6154) );
  INV_X1 U273 ( .A(n5120), .ZN(n6194) );
  INV_X1 U274 ( .A(n5119), .ZN(n6186) );
  INV_X1 U275 ( .A(n5139), .ZN(n6127) );
  INV_X1 U276 ( .A(n5138), .ZN(n6119) );
  INV_X1 U277 ( .A(n5144), .ZN(n6100) );
  INV_X1 U278 ( .A(n5143), .ZN(n6092) );
  BUF_X1 U279 ( .A(n1684), .Z(n6753) );
  BUF_X1 U280 ( .A(n1684), .Z(n6752) );
  BUF_X1 U281 ( .A(n1684), .Z(n6751) );
  BUF_X1 U282 ( .A(n1684), .Z(n6750) );
  BUF_X1 U283 ( .A(n1684), .Z(n6749) );
  BUF_X1 U284 ( .A(n1684), .Z(n6748) );
  INV_X1 U285 ( .A(n5115), .ZN(n6226) );
  INV_X1 U286 ( .A(n5114), .ZN(n6218) );
  INV_X1 U287 ( .A(n2896), .ZN(n6577) );
  INV_X1 U288 ( .A(n2896), .ZN(n6576) );
  INV_X1 U289 ( .A(n2861), .ZN(n6586) );
  INV_X1 U290 ( .A(n2861), .ZN(n6585) );
  INV_X1 U291 ( .A(n2619), .ZN(n6646) );
  INV_X1 U292 ( .A(n2619), .ZN(n6645) );
  INV_X1 U293 ( .A(n2584), .ZN(n6655) );
  INV_X1 U294 ( .A(n2584), .ZN(n6654) );
  INV_X1 U295 ( .A(n1897), .ZN(n6714) );
  INV_X1 U296 ( .A(n1897), .ZN(n6713) );
  INV_X1 U297 ( .A(n1862), .ZN(n6723) );
  INV_X1 U298 ( .A(n1862), .ZN(n6722) );
  INV_X1 U299 ( .A(n4320), .ZN(n6509) );
  INV_X1 U300 ( .A(n4320), .ZN(n6510) );
  INV_X1 U301 ( .A(n4285), .ZN(n6517) );
  INV_X1 U302 ( .A(n4285), .ZN(n6518) );
  INV_X1 U303 ( .A(n4183), .ZN(n6542) );
  INV_X1 U304 ( .A(n4183), .ZN(n6543) );
  INV_X1 U305 ( .A(n4148), .ZN(n6550) );
  INV_X1 U306 ( .A(n4148), .ZN(n6551) );
  INV_X1 U307 ( .A(n2756), .ZN(n6611) );
  INV_X1 U308 ( .A(n2756), .ZN(n6612) );
  INV_X1 U309 ( .A(n2721), .ZN(n6619) );
  INV_X1 U310 ( .A(n2721), .ZN(n6620) );
  INV_X1 U311 ( .A(n2032), .ZN(n6681) );
  INV_X1 U312 ( .A(n2032), .ZN(n6682) );
  INV_X1 U313 ( .A(n1997), .ZN(n6690) );
  INV_X1 U314 ( .A(n1997), .ZN(n6691) );
  BUF_X1 U315 ( .A(n1684), .Z(n6754) );
  INV_X1 U316 ( .A(n6731), .ZN(n1823) );
  INV_X1 U317 ( .A(n6733), .ZN(n1788) );
  BUF_X1 U318 ( .A(n6173), .Z(n6174) );
  BUF_X1 U319 ( .A(n6173), .Z(n6175) );
  BUF_X1 U320 ( .A(n6265), .Z(n6266) );
  BUF_X1 U321 ( .A(n6265), .Z(n6267) );
  INV_X1 U322 ( .A(n4391), .ZN(n6492) );
  INV_X1 U323 ( .A(n4391), .ZN(n6491) );
  INV_X1 U324 ( .A(n4357), .ZN(n6501) );
  INV_X1 U325 ( .A(n4357), .ZN(n6500) );
  INV_X1 U326 ( .A(n2973), .ZN(n6559) );
  INV_X1 U327 ( .A(n2973), .ZN(n6558) );
  INV_X1 U328 ( .A(n2930), .ZN(n6568) );
  INV_X1 U329 ( .A(n2930), .ZN(n6567) );
  INV_X1 U330 ( .A(n2687), .ZN(n6628) );
  INV_X1 U331 ( .A(n2687), .ZN(n6627) );
  INV_X1 U332 ( .A(n2653), .ZN(n6637) );
  INV_X1 U333 ( .A(n2653), .ZN(n6636) );
  INV_X1 U334 ( .A(n4251), .ZN(n6525) );
  INV_X1 U335 ( .A(n4251), .ZN(n6526) );
  INV_X1 U336 ( .A(n4217), .ZN(n6533) );
  INV_X1 U337 ( .A(n2824), .ZN(n6594) );
  INV_X1 U338 ( .A(n2824), .ZN(n6595) );
  INV_X1 U339 ( .A(n2790), .ZN(n6602) );
  INV_X1 U340 ( .A(n2100), .ZN(n6663) );
  INV_X1 U341 ( .A(n2100), .ZN(n6664) );
  INV_X1 U342 ( .A(n2066), .ZN(n6672) );
  INV_X1 U343 ( .A(n2066), .ZN(n6673) );
  BUF_X1 U344 ( .A(n6699), .Z(n6700) );
  BUF_X1 U345 ( .A(n6706), .Z(n6707) );
  BUF_X1 U346 ( .A(n6699), .Z(n6701) );
  BUF_X1 U347 ( .A(n6699), .Z(n6702) );
  BUF_X1 U348 ( .A(n6706), .Z(n6708) );
  BUF_X1 U349 ( .A(n6706), .Z(n6709) );
  BUF_X1 U350 ( .A(n6173), .Z(n6176) );
  BUF_X1 U351 ( .A(n5128), .Z(n6177) );
  BUF_X1 U352 ( .A(n5128), .Z(n6178) );
  BUF_X1 U353 ( .A(n5128), .Z(n6179) );
  BUF_X1 U354 ( .A(n6265), .Z(n6268) );
  BUF_X1 U355 ( .A(n5104), .Z(n6269) );
  BUF_X1 U356 ( .A(n5104), .Z(n6270) );
  BUF_X1 U357 ( .A(n5104), .Z(n6271) );
  INV_X1 U358 ( .A(add_rd2[2]), .ZN(n5080) );
  INV_X1 U359 ( .A(add_rd2[1]), .ZN(n5083) );
  BUF_X1 U360 ( .A(n1965), .Z(n6703) );
  BUF_X1 U361 ( .A(n1965), .Z(n6704) );
  BUF_X1 U362 ( .A(n1965), .Z(n6705) );
  BUF_X1 U363 ( .A(n1931), .Z(n6710) );
  BUF_X1 U364 ( .A(n1931), .Z(n6711) );
  BUF_X1 U365 ( .A(n1931), .Z(n6712) );
  BUF_X1 U366 ( .A(reset), .Z(n6763) );
  BUF_X1 U367 ( .A(reset), .Z(n6764) );
  BUF_X1 U368 ( .A(reset), .Z(n6765) );
  INV_X1 U369 ( .A(datain[0]), .ZN(n1748) );
  INV_X1 U370 ( .A(datain[1]), .ZN(n1746) );
  INV_X1 U371 ( .A(datain[2]), .ZN(n1744) );
  INV_X1 U372 ( .A(datain[3]), .ZN(n1742) );
  INV_X1 U373 ( .A(datain[4]), .ZN(n1740) );
  INV_X1 U374 ( .A(datain[5]), .ZN(n1738) );
  INV_X1 U375 ( .A(datain[6]), .ZN(n1736) );
  INV_X1 U376 ( .A(datain[7]), .ZN(n1734) );
  INV_X1 U377 ( .A(datain[8]), .ZN(n1732) );
  INV_X1 U378 ( .A(datain[9]), .ZN(n1730) );
  INV_X1 U379 ( .A(datain[10]), .ZN(n1728) );
  INV_X1 U380 ( .A(datain[11]), .ZN(n1726) );
  INV_X1 U381 ( .A(datain[12]), .ZN(n1724) );
  INV_X1 U382 ( .A(datain[13]), .ZN(n1722) );
  INV_X1 U383 ( .A(datain[14]), .ZN(n1720) );
  INV_X1 U384 ( .A(datain[15]), .ZN(n1718) );
  INV_X1 U385 ( .A(datain[16]), .ZN(n1716) );
  INV_X1 U386 ( .A(datain[17]), .ZN(n1714) );
  INV_X1 U387 ( .A(datain[18]), .ZN(n1712) );
  INV_X1 U388 ( .A(datain[19]), .ZN(n1710) );
  INV_X1 U389 ( .A(datain[20]), .ZN(n1708) );
  INV_X1 U390 ( .A(datain[21]), .ZN(n1706) );
  INV_X1 U391 ( .A(datain[22]), .ZN(n1704) );
  INV_X1 U392 ( .A(datain[23]), .ZN(n1702) );
  INV_X1 U393 ( .A(datain[24]), .ZN(n1700) );
  INV_X1 U394 ( .A(datain[25]), .ZN(n1698) );
  INV_X1 U395 ( .A(datain[26]), .ZN(n1696) );
  INV_X1 U396 ( .A(datain[27]), .ZN(n1694) );
  INV_X1 U397 ( .A(datain[28]), .ZN(n1692) );
  INV_X1 U398 ( .A(datain[29]), .ZN(n1690) );
  INV_X1 U399 ( .A(datain[30]), .ZN(n1688) );
  INV_X1 U400 ( .A(datain[31]), .ZN(n1685) );
  NOR3_X1 U401 ( .A1(n5744), .A2(n5748), .A3(n5745), .ZN(n5737) );
  NOR2_X1 U402 ( .A1(n5751), .A2(n5749), .ZN(n5738) );
  NAND2_X1 U403 ( .A1(n5736), .A2(n5729), .ZN(n6180) );
  NAND2_X1 U404 ( .A1(n5736), .A2(n5729), .ZN(n6181) );
  NAND2_X1 U405 ( .A1(n1856), .A2(n1751), .ZN(n6732) );
  NAND2_X1 U406 ( .A1(n1856), .A2(n1751), .ZN(n1822) );
  NAND2_X1 U407 ( .A1(n1821), .A2(n1751), .ZN(n6734) );
  NAND2_X1 U408 ( .A1(n1821), .A2(n1751), .ZN(n1787) );
  NAND2_X1 U409 ( .A1(n5724), .A2(n5725), .ZN(n6272) );
  NAND2_X1 U410 ( .A1(n5724), .A2(n5725), .ZN(n6273) );
  NAND2_X1 U411 ( .A1(n1856), .A2(n1751), .ZN(n6731) );
  NAND2_X1 U412 ( .A1(n1821), .A2(n1751), .ZN(n6733) );
  NAND2_X1 U413 ( .A1(n5736), .A2(n5729), .ZN(n5129) );
  NAND2_X1 U414 ( .A1(n5724), .A2(n5725), .ZN(n5105) );
  AND2_X1 U415 ( .A1(n5727), .A2(n5726), .ZN(n6261) );
  AND2_X1 U416 ( .A1(n5727), .A2(n5726), .ZN(n6262) );
  AND2_X1 U417 ( .A1(n5727), .A2(n5725), .ZN(n6263) );
  AND2_X1 U418 ( .A1(n5727), .A2(n5725), .ZN(n6264) );
  AND2_X1 U419 ( .A1(n5735), .A2(n5738), .ZN(n6184) );
  AND2_X1 U420 ( .A1(n5735), .A2(n5738), .ZN(n6185) );
  AND2_X1 U421 ( .A1(n5727), .A2(n5726), .ZN(n5101) );
  AND2_X1 U422 ( .A1(n5727), .A2(n5725), .ZN(n5102) );
  AND2_X1 U423 ( .A1(n5735), .A2(n5738), .ZN(n5117) );
  AND3_X1 U424 ( .A1(n1857), .A2(n1858), .A3(n1859), .ZN(n1751) );
  NAND2_X1 U425 ( .A1(n5725), .A2(n5736), .ZN(n5133) );
  NAND2_X1 U426 ( .A1(n5724), .A2(n5729), .ZN(n5110) );
  NAND2_X1 U427 ( .A1(n5724), .A2(n5730), .ZN(n5109) );
  NAND2_X1 U428 ( .A1(n5726), .A2(n5736), .ZN(n5134) );
  NAND2_X1 U429 ( .A1(n5724), .A2(n5726), .ZN(n6265) );
  NAND2_X1 U430 ( .A1(n5724), .A2(n5726), .ZN(n5104) );
  NAND2_X1 U431 ( .A1(n1750), .A2(n1751), .ZN(n1684) );
  NAND2_X1 U432 ( .A1(n5737), .A2(n5736), .ZN(n5119) );
  NAND2_X1 U433 ( .A1(n5737), .A2(n5724), .ZN(n5138) );
  NAND2_X1 U434 ( .A1(n5735), .A2(n5736), .ZN(n5120) );
  NAND2_X1 U435 ( .A1(n5735), .A2(n5724), .ZN(n5139) );
  INV_X1 U436 ( .A(n5718), .ZN(n5752) );
  INV_X1 U437 ( .A(n5050), .ZN(n5084) );
  NAND2_X1 U438 ( .A1(n5732), .A2(n5736), .ZN(n5144) );
  NAND2_X1 U439 ( .A1(n5733), .A2(n5736), .ZN(n5143) );
  OAI22_X1 U440 ( .A1(n1748), .A2(n6516), .B1(n5988), .B2(n4246), .ZN(n3179)
         );
  OAI22_X1 U441 ( .A1(n1746), .A2(n6511), .B1(n5988), .B2(n4247), .ZN(n3180)
         );
  OAI22_X1 U442 ( .A1(n1744), .A2(n6511), .B1(n5988), .B2(n4248), .ZN(n3181)
         );
  OAI22_X1 U443 ( .A1(n1742), .A2(n6514), .B1(n5988), .B2(n4249), .ZN(n3182)
         );
  OAI22_X1 U444 ( .A1(n1740), .A2(n6511), .B1(n5988), .B2(n4250), .ZN(n3183)
         );
  OAI22_X1 U445 ( .A1(n1738), .A2(n6512), .B1(n5988), .B2(n4253), .ZN(n3184)
         );
  OAI22_X1 U446 ( .A1(n1736), .A2(n6513), .B1(n5988), .B2(n4254), .ZN(n3185)
         );
  OAI22_X1 U447 ( .A1(n1734), .A2(n6513), .B1(n5988), .B2(n4255), .ZN(n3186)
         );
  OAI22_X1 U448 ( .A1(n1732), .A2(n6514), .B1(n5988), .B2(n4256), .ZN(n3187)
         );
  OAI22_X1 U449 ( .A1(n1730), .A2(n6514), .B1(n5988), .B2(n4257), .ZN(n3188)
         );
  OAI22_X1 U450 ( .A1(n1728), .A2(n6515), .B1(n5988), .B2(n4258), .ZN(n3189)
         );
  OAI22_X1 U451 ( .A1(n1726), .A2(n6511), .B1(n5988), .B2(n4259), .ZN(n3190)
         );
  OAI22_X1 U452 ( .A1(n1724), .A2(n6513), .B1(n5989), .B2(n4260), .ZN(n3191)
         );
  OAI22_X1 U453 ( .A1(n1722), .A2(n6513), .B1(n5989), .B2(n4261), .ZN(n3192)
         );
  OAI22_X1 U454 ( .A1(n1720), .A2(n6515), .B1(n5989), .B2(n4262), .ZN(n3193)
         );
  OAI22_X1 U455 ( .A1(n1718), .A2(n6514), .B1(n5989), .B2(n4263), .ZN(n3194)
         );
  OAI22_X1 U456 ( .A1(n1716), .A2(n6515), .B1(n5989), .B2(n4264), .ZN(n3195)
         );
  OAI22_X1 U457 ( .A1(n1714), .A2(n6511), .B1(n5989), .B2(n4265), .ZN(n3196)
         );
  OAI22_X1 U458 ( .A1(n1712), .A2(n6515), .B1(n5989), .B2(n4266), .ZN(n3197)
         );
  OAI22_X1 U459 ( .A1(n1710), .A2(n6511), .B1(n5989), .B2(n4267), .ZN(n3198)
         );
  OAI22_X1 U460 ( .A1(n1708), .A2(n6515), .B1(n5989), .B2(n4268), .ZN(n3199)
         );
  OAI22_X1 U461 ( .A1(n1706), .A2(n6516), .B1(n5989), .B2(n4269), .ZN(n3200)
         );
  OAI22_X1 U462 ( .A1(n1704), .A2(n6513), .B1(n5989), .B2(n4270), .ZN(n3201)
         );
  OAI22_X1 U463 ( .A1(n1702), .A2(n6514), .B1(n5989), .B2(n4271), .ZN(n3202)
         );
  OAI22_X1 U464 ( .A1(n1748), .A2(n6522), .B1(n5991), .B2(n5944), .ZN(n3211)
         );
  OAI22_X1 U465 ( .A1(n1746), .A2(n6523), .B1(n5991), .B2(n5945), .ZN(n3212)
         );
  OAI22_X1 U466 ( .A1(n1744), .A2(n6524), .B1(n5991), .B2(n5946), .ZN(n3213)
         );
  OAI22_X1 U467 ( .A1(n1742), .A2(n6521), .B1(n5991), .B2(n5947), .ZN(n3214)
         );
  OAI22_X1 U468 ( .A1(n1740), .A2(n6522), .B1(n5991), .B2(n5948), .ZN(n3215)
         );
  OAI22_X1 U469 ( .A1(n1738), .A2(n6519), .B1(n5991), .B2(n5949), .ZN(n3216)
         );
  OAI22_X1 U470 ( .A1(n1736), .A2(n6520), .B1(n5991), .B2(n5950), .ZN(n3217)
         );
  OAI22_X1 U471 ( .A1(n1734), .A2(n6520), .B1(n5991), .B2(n5951), .ZN(n3218)
         );
  OAI22_X1 U472 ( .A1(n1732), .A2(n6524), .B1(n5991), .B2(n5952), .ZN(n3219)
         );
  OAI22_X1 U473 ( .A1(n1730), .A2(n6521), .B1(n5991), .B2(n5953), .ZN(n3220)
         );
  OAI22_X1 U474 ( .A1(n1728), .A2(n6522), .B1(n5991), .B2(n5954), .ZN(n3221)
         );
  OAI22_X1 U475 ( .A1(n1726), .A2(n6523), .B1(n5991), .B2(n5955), .ZN(n3222)
         );
  OAI22_X1 U476 ( .A1(n1724), .A2(n6520), .B1(n5992), .B2(n5956), .ZN(n3223)
         );
  OAI22_X1 U477 ( .A1(n1722), .A2(n6520), .B1(n5992), .B2(n5957), .ZN(n3224)
         );
  OAI22_X1 U478 ( .A1(n1720), .A2(n6521), .B1(n5992), .B2(n5958), .ZN(n3225)
         );
  OAI22_X1 U479 ( .A1(n1718), .A2(n6521), .B1(n5992), .B2(n5959), .ZN(n3226)
         );
  OAI22_X1 U480 ( .A1(n1716), .A2(n6522), .B1(n5992), .B2(n5960), .ZN(n3227)
         );
  OAI22_X1 U481 ( .A1(n1714), .A2(n6523), .B1(n5992), .B2(n5961), .ZN(n3228)
         );
  OAI22_X1 U482 ( .A1(n1712), .A2(n6523), .B1(n5992), .B2(n5962), .ZN(n3229)
         );
  OAI22_X1 U483 ( .A1(n1710), .A2(n6522), .B1(n5992), .B2(n5963), .ZN(n3230)
         );
  OAI22_X1 U484 ( .A1(n1708), .A2(n6522), .B1(n5992), .B2(n5964), .ZN(n3231)
         );
  OAI22_X1 U485 ( .A1(n1706), .A2(n6523), .B1(n5992), .B2(n5965), .ZN(n3232)
         );
  OAI22_X1 U486 ( .A1(n1704), .A2(n6520), .B1(n5992), .B2(n5966), .ZN(n3233)
         );
  OAI22_X1 U487 ( .A1(n1702), .A2(n6524), .B1(n5992), .B2(n5967), .ZN(n3234)
         );
  OAI22_X1 U488 ( .A1(n1748), .A2(n6532), .B1(n5994), .B2(n2852), .ZN(n3243)
         );
  OAI22_X1 U489 ( .A1(n1746), .A2(n6527), .B1(n5994), .B2(n2854), .ZN(n3244)
         );
  OAI22_X1 U490 ( .A1(n1744), .A2(n6527), .B1(n5994), .B2(n2856), .ZN(n3245)
         );
  OAI22_X1 U491 ( .A1(n1742), .A2(n6530), .B1(n5994), .B2(n2860), .ZN(n3246)
         );
  OAI22_X1 U492 ( .A1(n1740), .A2(n6527), .B1(n5994), .B2(n2929), .ZN(n3247)
         );
  OAI22_X1 U493 ( .A1(n1738), .A2(n6528), .B1(n5994), .B2(n4150), .ZN(n3248)
         );
  OAI22_X1 U494 ( .A1(n1736), .A2(n6529), .B1(n5994), .B2(n4152), .ZN(n3249)
         );
  OAI22_X1 U495 ( .A1(n1734), .A2(n6529), .B1(n5994), .B2(n4154), .ZN(n3250)
         );
  OAI22_X1 U496 ( .A1(n1732), .A2(n6530), .B1(n5994), .B2(n4156), .ZN(n3251)
         );
  OAI22_X1 U497 ( .A1(n1730), .A2(n6530), .B1(n5994), .B2(n4158), .ZN(n3252)
         );
  OAI22_X1 U498 ( .A1(n1728), .A2(n6531), .B1(n5994), .B2(n4160), .ZN(n3253)
         );
  OAI22_X1 U499 ( .A1(n1726), .A2(n6527), .B1(n5994), .B2(n4162), .ZN(n3254)
         );
  OAI22_X1 U500 ( .A1(n1724), .A2(n6529), .B1(n5995), .B2(n4164), .ZN(n3255)
         );
  OAI22_X1 U501 ( .A1(n1722), .A2(n6529), .B1(n5995), .B2(n4166), .ZN(n3256)
         );
  OAI22_X1 U502 ( .A1(n1720), .A2(n6531), .B1(n5995), .B2(n4168), .ZN(n3257)
         );
  OAI22_X1 U503 ( .A1(n1718), .A2(n6530), .B1(n5995), .B2(n4170), .ZN(n3258)
         );
  OAI22_X1 U504 ( .A1(n1716), .A2(n6531), .B1(n5995), .B2(n4172), .ZN(n3259)
         );
  OAI22_X1 U505 ( .A1(n1714), .A2(n6527), .B1(n5995), .B2(n4174), .ZN(n3260)
         );
  OAI22_X1 U506 ( .A1(n1712), .A2(n6531), .B1(n5995), .B2(n4176), .ZN(n3261)
         );
  OAI22_X1 U507 ( .A1(n1710), .A2(n6527), .B1(n5995), .B2(n4178), .ZN(n3262)
         );
  OAI22_X1 U508 ( .A1(n1708), .A2(n6532), .B1(n5995), .B2(n4199), .ZN(n3263)
         );
  OAI22_X1 U509 ( .A1(n1706), .A2(n6531), .B1(n5995), .B2(n4200), .ZN(n3264)
         );
  OAI22_X1 U510 ( .A1(n1704), .A2(n6529), .B1(n5995), .B2(n4201), .ZN(n3265)
         );
  OAI22_X1 U511 ( .A1(n1702), .A2(n6530), .B1(n5995), .B2(n4203), .ZN(n3266)
         );
  OAI22_X1 U512 ( .A1(n1748), .A2(n6534), .B1(n5997), .B2(n5842), .ZN(n3275)
         );
  OAI22_X1 U513 ( .A1(n1746), .A2(n6535), .B1(n5997), .B2(n5844), .ZN(n3276)
         );
  OAI22_X1 U514 ( .A1(n1744), .A2(n6541), .B1(n5997), .B2(n5846), .ZN(n3277)
         );
  OAI22_X1 U515 ( .A1(n1742), .A2(n6536), .B1(n5997), .B2(n5848), .ZN(n3278)
         );
  OAI22_X1 U516 ( .A1(n1740), .A2(n6537), .B1(n5997), .B2(n5850), .ZN(n3279)
         );
  OAI22_X1 U517 ( .A1(n1738), .A2(n6539), .B1(n5997), .B2(n5852), .ZN(n3280)
         );
  OAI22_X1 U518 ( .A1(n1736), .A2(n6535), .B1(n5997), .B2(n5854), .ZN(n3281)
         );
  OAI22_X1 U519 ( .A1(n1734), .A2(n6536), .B1(n5997), .B2(n5856), .ZN(n3282)
         );
  OAI22_X1 U520 ( .A1(n1732), .A2(n6537), .B1(n5997), .B2(n5858), .ZN(n3283)
         );
  OAI22_X1 U521 ( .A1(n1730), .A2(n6540), .B1(n5997), .B2(n5860), .ZN(n3284)
         );
  OAI22_X1 U522 ( .A1(n1728), .A2(n6538), .B1(n5997), .B2(n5862), .ZN(n3285)
         );
  OAI22_X1 U523 ( .A1(n1726), .A2(n6539), .B1(n5997), .B2(n5864), .ZN(n3286)
         );
  OAI22_X1 U524 ( .A1(n1724), .A2(n6536), .B1(n5998), .B2(n5866), .ZN(n3287)
         );
  OAI22_X1 U525 ( .A1(n1722), .A2(n6537), .B1(n5998), .B2(n5868), .ZN(n3288)
         );
  OAI22_X1 U526 ( .A1(n1720), .A2(n6541), .B1(n5998), .B2(n5870), .ZN(n3289)
         );
  OAI22_X1 U527 ( .A1(n1718), .A2(n6534), .B1(n5998), .B2(n5872), .ZN(n3290)
         );
  OAI22_X1 U528 ( .A1(n1716), .A2(n6538), .B1(n5998), .B2(n5874), .ZN(n3291)
         );
  OAI22_X1 U529 ( .A1(n1714), .A2(n6539), .B1(n5998), .B2(n5876), .ZN(n3292)
         );
  OAI22_X1 U530 ( .A1(n1712), .A2(n6540), .B1(n5998), .B2(n5878), .ZN(n3293)
         );
  OAI22_X1 U531 ( .A1(n1710), .A2(n6537), .B1(n5998), .B2(n5880), .ZN(n3294)
         );
  OAI22_X1 U532 ( .A1(n1708), .A2(n6540), .B1(n5998), .B2(n5898), .ZN(n3295)
         );
  OAI22_X1 U533 ( .A1(n1706), .A2(n6539), .B1(n5998), .B2(n5899), .ZN(n3296)
         );
  OAI22_X1 U534 ( .A1(n1704), .A2(n6535), .B1(n5998), .B2(n5900), .ZN(n3297)
         );
  OAI22_X1 U535 ( .A1(n1702), .A2(n6541), .B1(n5998), .B2(n5902), .ZN(n3298)
         );
  OAI22_X1 U536 ( .A1(n1748), .A2(n6549), .B1(n6000), .B2(n4220), .ZN(n3307)
         );
  OAI22_X1 U537 ( .A1(n1746), .A2(n6544), .B1(n6000), .B2(n4221), .ZN(n3308)
         );
  OAI22_X1 U538 ( .A1(n1744), .A2(n6544), .B1(n6000), .B2(n4222), .ZN(n3309)
         );
  OAI22_X1 U539 ( .A1(n1742), .A2(n6547), .B1(n6000), .B2(n4223), .ZN(n3310)
         );
  OAI22_X1 U540 ( .A1(n1740), .A2(n6544), .B1(n6000), .B2(n4224), .ZN(n3311)
         );
  OAI22_X1 U541 ( .A1(n1738), .A2(n6545), .B1(n6000), .B2(n4225), .ZN(n3312)
         );
  OAI22_X1 U542 ( .A1(n1736), .A2(n6546), .B1(n6000), .B2(n4226), .ZN(n3313)
         );
  OAI22_X1 U543 ( .A1(n1734), .A2(n6546), .B1(n6000), .B2(n4227), .ZN(n3314)
         );
  OAI22_X1 U544 ( .A1(n1732), .A2(n6547), .B1(n6000), .B2(n4228), .ZN(n3315)
         );
  OAI22_X1 U545 ( .A1(n1730), .A2(n6547), .B1(n6000), .B2(n4229), .ZN(n3316)
         );
  OAI22_X1 U546 ( .A1(n1728), .A2(n6548), .B1(n6000), .B2(n4230), .ZN(n3317)
         );
  OAI22_X1 U547 ( .A1(n1726), .A2(n6544), .B1(n6000), .B2(n4231), .ZN(n3318)
         );
  OAI22_X1 U548 ( .A1(n1724), .A2(n6546), .B1(n6001), .B2(n4232), .ZN(n3319)
         );
  OAI22_X1 U549 ( .A1(n1722), .A2(n6546), .B1(n6001), .B2(n4233), .ZN(n3320)
         );
  OAI22_X1 U550 ( .A1(n1720), .A2(n6548), .B1(n6001), .B2(n4234), .ZN(n3321)
         );
  OAI22_X1 U551 ( .A1(n1718), .A2(n6547), .B1(n6001), .B2(n4235), .ZN(n3322)
         );
  OAI22_X1 U552 ( .A1(n1716), .A2(n6548), .B1(n6001), .B2(n4236), .ZN(n3323)
         );
  OAI22_X1 U553 ( .A1(n1714), .A2(n6544), .B1(n6001), .B2(n4237), .ZN(n3324)
         );
  OAI22_X1 U554 ( .A1(n1712), .A2(n6548), .B1(n6001), .B2(n4238), .ZN(n3325)
         );
  OAI22_X1 U555 ( .A1(n1710), .A2(n6544), .B1(n6001), .B2(n4239), .ZN(n3326)
         );
  OAI22_X1 U556 ( .A1(n1708), .A2(n6548), .B1(n6001), .B2(n4240), .ZN(n3327)
         );
  OAI22_X1 U557 ( .A1(n1706), .A2(n6549), .B1(n6001), .B2(n4241), .ZN(n3328)
         );
  OAI22_X1 U558 ( .A1(n1704), .A2(n6546), .B1(n6001), .B2(n4280), .ZN(n3329)
         );
  OAI22_X1 U559 ( .A1(n1702), .A2(n6547), .B1(n6001), .B2(n4281), .ZN(n3330)
         );
  OAI22_X1 U560 ( .A1(n1748), .A2(n6555), .B1(n6003), .B2(n5918), .ZN(n3339)
         );
  OAI22_X1 U561 ( .A1(n1746), .A2(n6556), .B1(n6003), .B2(n5919), .ZN(n3340)
         );
  OAI22_X1 U562 ( .A1(n1744), .A2(n6557), .B1(n6003), .B2(n5920), .ZN(n3341)
         );
  OAI22_X1 U563 ( .A1(n1742), .A2(n6554), .B1(n6003), .B2(n5921), .ZN(n3342)
         );
  OAI22_X1 U564 ( .A1(n1740), .A2(n6555), .B1(n6003), .B2(n5922), .ZN(n3343)
         );
  OAI22_X1 U565 ( .A1(n1738), .A2(n6552), .B1(n6003), .B2(n5923), .ZN(n3344)
         );
  OAI22_X1 U566 ( .A1(n1736), .A2(n6553), .B1(n6003), .B2(n5924), .ZN(n3345)
         );
  OAI22_X1 U567 ( .A1(n1734), .A2(n6553), .B1(n6003), .B2(n5925), .ZN(n3346)
         );
  OAI22_X1 U568 ( .A1(n1732), .A2(n6557), .B1(n6003), .B2(n5926), .ZN(n3347)
         );
  OAI22_X1 U569 ( .A1(n1730), .A2(n6554), .B1(n6003), .B2(n5927), .ZN(n3348)
         );
  OAI22_X1 U570 ( .A1(n1728), .A2(n6555), .B1(n6003), .B2(n5928), .ZN(n3349)
         );
  OAI22_X1 U571 ( .A1(n1726), .A2(n6556), .B1(n6003), .B2(n5929), .ZN(n3350)
         );
  OAI22_X1 U572 ( .A1(n1724), .A2(n6553), .B1(n6004), .B2(n5930), .ZN(n3351)
         );
  OAI22_X1 U573 ( .A1(n1722), .A2(n6553), .B1(n6004), .B2(n5931), .ZN(n3352)
         );
  OAI22_X1 U574 ( .A1(n1720), .A2(n6554), .B1(n6004), .B2(n5932), .ZN(n3353)
         );
  OAI22_X1 U575 ( .A1(n1718), .A2(n6554), .B1(n6004), .B2(n5933), .ZN(n3354)
         );
  OAI22_X1 U576 ( .A1(n1716), .A2(n6555), .B1(n6004), .B2(n5934), .ZN(n3355)
         );
  OAI22_X1 U577 ( .A1(n1714), .A2(n6556), .B1(n6004), .B2(n5935), .ZN(n3356)
         );
  OAI22_X1 U578 ( .A1(n1712), .A2(n6556), .B1(n6004), .B2(n5936), .ZN(n3357)
         );
  OAI22_X1 U579 ( .A1(n1710), .A2(n6555), .B1(n6004), .B2(n5937), .ZN(n3358)
         );
  OAI22_X1 U580 ( .A1(n1708), .A2(n6555), .B1(n6004), .B2(n5938), .ZN(n3359)
         );
  OAI22_X1 U581 ( .A1(n1706), .A2(n6556), .B1(n6004), .B2(n5939), .ZN(n3360)
         );
  OAI22_X1 U582 ( .A1(n1704), .A2(n6553), .B1(n6004), .B2(n5976), .ZN(n3361)
         );
  OAI22_X1 U583 ( .A1(n1702), .A2(n6557), .B1(n6004), .B2(n5977), .ZN(n3362)
         );
  OAI22_X1 U584 ( .A1(n1748), .A2(n6601), .B1(n6018), .B2(n2853), .ZN(n3499)
         );
  OAI22_X1 U585 ( .A1(n1746), .A2(n6596), .B1(n6018), .B2(n2855), .ZN(n3500)
         );
  OAI22_X1 U586 ( .A1(n1744), .A2(n6596), .B1(n6018), .B2(n2857), .ZN(n3501)
         );
  OAI22_X1 U587 ( .A1(n1742), .A2(n6599), .B1(n6018), .B2(n2895), .ZN(n3502)
         );
  OAI22_X1 U588 ( .A1(n1740), .A2(n6596), .B1(n6018), .B2(n2971), .ZN(n3503)
         );
  OAI22_X1 U589 ( .A1(n1738), .A2(n6597), .B1(n6018), .B2(n4151), .ZN(n3504)
         );
  OAI22_X1 U590 ( .A1(n1736), .A2(n6598), .B1(n6018), .B2(n4153), .ZN(n3505)
         );
  OAI22_X1 U591 ( .A1(n1734), .A2(n6598), .B1(n6018), .B2(n4155), .ZN(n3506)
         );
  OAI22_X1 U592 ( .A1(n1732), .A2(n6599), .B1(n6018), .B2(n4157), .ZN(n3507)
         );
  OAI22_X1 U593 ( .A1(n1730), .A2(n6599), .B1(n6018), .B2(n4159), .ZN(n3508)
         );
  OAI22_X1 U594 ( .A1(n1728), .A2(n6600), .B1(n6018), .B2(n4161), .ZN(n3509)
         );
  OAI22_X1 U595 ( .A1(n1726), .A2(n6596), .B1(n6018), .B2(n4163), .ZN(n3510)
         );
  OAI22_X1 U596 ( .A1(n1724), .A2(n6598), .B1(n6019), .B2(n4165), .ZN(n3511)
         );
  OAI22_X1 U597 ( .A1(n1722), .A2(n6598), .B1(n6019), .B2(n4167), .ZN(n3512)
         );
  OAI22_X1 U598 ( .A1(n1720), .A2(n6600), .B1(n6019), .B2(n4169), .ZN(n3513)
         );
  OAI22_X1 U599 ( .A1(n1718), .A2(n6599), .B1(n6019), .B2(n4171), .ZN(n3514)
         );
  OAI22_X1 U600 ( .A1(n1716), .A2(n6600), .B1(n6019), .B2(n4173), .ZN(n3515)
         );
  OAI22_X1 U601 ( .A1(n1714), .A2(n6596), .B1(n6019), .B2(n4175), .ZN(n3516)
         );
  OAI22_X1 U602 ( .A1(n1712), .A2(n6600), .B1(n6019), .B2(n4177), .ZN(n3517)
         );
  OAI22_X1 U603 ( .A1(n1710), .A2(n6596), .B1(n6019), .B2(n4179), .ZN(n3518)
         );
  OAI22_X1 U604 ( .A1(n1708), .A2(n6601), .B1(n6019), .B2(n4180), .ZN(n3519)
         );
  OAI22_X1 U605 ( .A1(n1706), .A2(n6600), .B1(n6019), .B2(n4181), .ZN(n3520)
         );
  OAI22_X1 U606 ( .A1(n1704), .A2(n6598), .B1(n6019), .B2(n4185), .ZN(n3521)
         );
  OAI22_X1 U607 ( .A1(n1702), .A2(n6599), .B1(n6019), .B2(n4186), .ZN(n3522)
         );
  OAI22_X1 U608 ( .A1(n1748), .A2(n6603), .B1(n6021), .B2(n5843), .ZN(n3531)
         );
  OAI22_X1 U609 ( .A1(n1746), .A2(n6604), .B1(n6021), .B2(n5845), .ZN(n3532)
         );
  OAI22_X1 U610 ( .A1(n1744), .A2(n6610), .B1(n6021), .B2(n5847), .ZN(n3533)
         );
  OAI22_X1 U611 ( .A1(n1742), .A2(n6605), .B1(n6021), .B2(n5849), .ZN(n3534)
         );
  OAI22_X1 U612 ( .A1(n1740), .A2(n6606), .B1(n6021), .B2(n5851), .ZN(n3535)
         );
  OAI22_X1 U613 ( .A1(n1738), .A2(n6608), .B1(n6021), .B2(n5853), .ZN(n3536)
         );
  OAI22_X1 U614 ( .A1(n1736), .A2(n6604), .B1(n6021), .B2(n5855), .ZN(n3537)
         );
  OAI22_X1 U615 ( .A1(n1734), .A2(n6605), .B1(n6021), .B2(n5857), .ZN(n3538)
         );
  OAI22_X1 U616 ( .A1(n1732), .A2(n6606), .B1(n6021), .B2(n5859), .ZN(n3539)
         );
  OAI22_X1 U617 ( .A1(n1730), .A2(n6609), .B1(n6021), .B2(n5861), .ZN(n3540)
         );
  OAI22_X1 U618 ( .A1(n1728), .A2(n6607), .B1(n6021), .B2(n5863), .ZN(n3541)
         );
  OAI22_X1 U619 ( .A1(n1726), .A2(n6608), .B1(n6021), .B2(n5865), .ZN(n3542)
         );
  OAI22_X1 U620 ( .A1(n1724), .A2(n6605), .B1(n6022), .B2(n5867), .ZN(n3543)
         );
  OAI22_X1 U621 ( .A1(n1722), .A2(n6606), .B1(n6022), .B2(n5869), .ZN(n3544)
         );
  OAI22_X1 U622 ( .A1(n1720), .A2(n6610), .B1(n6022), .B2(n5871), .ZN(n3545)
         );
  OAI22_X1 U623 ( .A1(n1718), .A2(n6603), .B1(n6022), .B2(n5873), .ZN(n3546)
         );
  OAI22_X1 U624 ( .A1(n1716), .A2(n6607), .B1(n6022), .B2(n5875), .ZN(n3547)
         );
  OAI22_X1 U625 ( .A1(n1714), .A2(n6608), .B1(n6022), .B2(n5877), .ZN(n3548)
         );
  OAI22_X1 U626 ( .A1(n1712), .A2(n6609), .B1(n6022), .B2(n5879), .ZN(n3549)
         );
  OAI22_X1 U627 ( .A1(n1710), .A2(n6606), .B1(n6022), .B2(n5881), .ZN(n3550)
         );
  OAI22_X1 U628 ( .A1(n1708), .A2(n6609), .B1(n6022), .B2(n5882), .ZN(n3551)
         );
  OAI22_X1 U629 ( .A1(n1706), .A2(n6608), .B1(n6022), .B2(n5883), .ZN(n3552)
         );
  OAI22_X1 U630 ( .A1(n1704), .A2(n6604), .B1(n6022), .B2(n5884), .ZN(n3553)
         );
  OAI22_X1 U631 ( .A1(n1702), .A2(n6610), .B1(n6022), .B2(n5885), .ZN(n3554)
         );
  OAI22_X1 U632 ( .A1(n1748), .A2(n6618), .B1(n6024), .B2(n2793), .ZN(n3563)
         );
  OAI22_X1 U633 ( .A1(n1746), .A2(n6613), .B1(n6024), .B2(n2795), .ZN(n3564)
         );
  OAI22_X1 U634 ( .A1(n1744), .A2(n6613), .B1(n6024), .B2(n2797), .ZN(n3565)
         );
  OAI22_X1 U635 ( .A1(n1742), .A2(n6616), .B1(n6024), .B2(n2799), .ZN(n3566)
         );
  OAI22_X1 U636 ( .A1(n1740), .A2(n6613), .B1(n6024), .B2(n2801), .ZN(n3567)
         );
  OAI22_X1 U637 ( .A1(n1738), .A2(n6614), .B1(n6024), .B2(n2803), .ZN(n3568)
         );
  OAI22_X1 U638 ( .A1(n1736), .A2(n6615), .B1(n6024), .B2(n2805), .ZN(n3569)
         );
  OAI22_X1 U639 ( .A1(n1734), .A2(n6615), .B1(n6024), .B2(n2807), .ZN(n3570)
         );
  OAI22_X1 U640 ( .A1(n1732), .A2(n6616), .B1(n6024), .B2(n2809), .ZN(n3571)
         );
  OAI22_X1 U641 ( .A1(n1730), .A2(n6616), .B1(n6024), .B2(n2811), .ZN(n3572)
         );
  OAI22_X1 U642 ( .A1(n1728), .A2(n6617), .B1(n6024), .B2(n2813), .ZN(n3573)
         );
  OAI22_X1 U643 ( .A1(n1726), .A2(n6613), .B1(n6024), .B2(n2815), .ZN(n3574)
         );
  OAI22_X1 U644 ( .A1(n1724), .A2(n6615), .B1(n6025), .B2(n2817), .ZN(n3575)
         );
  OAI22_X1 U645 ( .A1(n1722), .A2(n6615), .B1(n6025), .B2(n2819), .ZN(n3576)
         );
  OAI22_X1 U646 ( .A1(n1720), .A2(n6617), .B1(n6025), .B2(n2821), .ZN(n3577)
         );
  OAI22_X1 U647 ( .A1(n1718), .A2(n6616), .B1(n6025), .B2(n2823), .ZN(n3578)
         );
  OAI22_X1 U648 ( .A1(n1716), .A2(n6617), .B1(n6025), .B2(n2827), .ZN(n3579)
         );
  OAI22_X1 U649 ( .A1(n1714), .A2(n6613), .B1(n6025), .B2(n2829), .ZN(n3580)
         );
  OAI22_X1 U650 ( .A1(n1712), .A2(n6617), .B1(n6025), .B2(n2831), .ZN(n3581)
         );
  OAI22_X1 U651 ( .A1(n1710), .A2(n6613), .B1(n6025), .B2(n2833), .ZN(n3582)
         );
  OAI22_X1 U652 ( .A1(n1708), .A2(n6617), .B1(n6025), .B2(n2835), .ZN(n3583)
         );
  OAI22_X1 U653 ( .A1(n1706), .A2(n6618), .B1(n6025), .B2(n2837), .ZN(n3584)
         );
  OAI22_X1 U654 ( .A1(n1704), .A2(n6615), .B1(n6025), .B2(n4213), .ZN(n3585)
         );
  OAI22_X1 U655 ( .A1(n1702), .A2(n6616), .B1(n6025), .B2(n4214), .ZN(n3586)
         );
  OAI22_X1 U656 ( .A1(n1748), .A2(n6624), .B1(n6027), .B2(n5785), .ZN(n3595)
         );
  OAI22_X1 U657 ( .A1(n1746), .A2(n6625), .B1(n6027), .B2(n5787), .ZN(n3596)
         );
  OAI22_X1 U658 ( .A1(n1744), .A2(n6626), .B1(n6027), .B2(n5789), .ZN(n3597)
         );
  OAI22_X1 U659 ( .A1(n1742), .A2(n6623), .B1(n6027), .B2(n5791), .ZN(n3598)
         );
  OAI22_X1 U660 ( .A1(n1740), .A2(n6624), .B1(n6027), .B2(n5793), .ZN(n3599)
         );
  OAI22_X1 U661 ( .A1(n1738), .A2(n6621), .B1(n6027), .B2(n5795), .ZN(n3600)
         );
  OAI22_X1 U662 ( .A1(n1736), .A2(n6622), .B1(n6027), .B2(n5797), .ZN(n3601)
         );
  OAI22_X1 U663 ( .A1(n1734), .A2(n6622), .B1(n6027), .B2(n5799), .ZN(n3602)
         );
  OAI22_X1 U664 ( .A1(n1732), .A2(n6626), .B1(n6027), .B2(n5801), .ZN(n3603)
         );
  OAI22_X1 U665 ( .A1(n1730), .A2(n6623), .B1(n6027), .B2(n5803), .ZN(n3604)
         );
  OAI22_X1 U666 ( .A1(n1728), .A2(n6624), .B1(n6027), .B2(n5805), .ZN(n3605)
         );
  OAI22_X1 U667 ( .A1(n1726), .A2(n6625), .B1(n6027), .B2(n5807), .ZN(n3606)
         );
  OAI22_X1 U668 ( .A1(n1724), .A2(n6622), .B1(n6028), .B2(n5809), .ZN(n3607)
         );
  OAI22_X1 U669 ( .A1(n1722), .A2(n6622), .B1(n6028), .B2(n5811), .ZN(n3608)
         );
  OAI22_X1 U670 ( .A1(n1720), .A2(n6623), .B1(n6028), .B2(n5813), .ZN(n3609)
         );
  OAI22_X1 U671 ( .A1(n1718), .A2(n6623), .B1(n6028), .B2(n5815), .ZN(n3610)
         );
  OAI22_X1 U672 ( .A1(n1716), .A2(n6624), .B1(n6028), .B2(n5817), .ZN(n3611)
         );
  OAI22_X1 U673 ( .A1(n1714), .A2(n6625), .B1(n6028), .B2(n5819), .ZN(n3612)
         );
  OAI22_X1 U674 ( .A1(n1712), .A2(n6625), .B1(n6028), .B2(n5821), .ZN(n3613)
         );
  OAI22_X1 U675 ( .A1(n1710), .A2(n6624), .B1(n6028), .B2(n5823), .ZN(n3614)
         );
  OAI22_X1 U676 ( .A1(n1708), .A2(n6624), .B1(n6028), .B2(n5825), .ZN(n3615)
         );
  OAI22_X1 U677 ( .A1(n1706), .A2(n6625), .B1(n6028), .B2(n5827), .ZN(n3616)
         );
  OAI22_X1 U678 ( .A1(n1704), .A2(n6622), .B1(n6028), .B2(n5912), .ZN(n3617)
         );
  OAI22_X1 U679 ( .A1(n1702), .A2(n6626), .B1(n6028), .B2(n5913), .ZN(n3618)
         );
  OAI22_X1 U680 ( .A1(n1748), .A2(n6666), .B1(n6042), .B2(n2732), .ZN(n3755)
         );
  OAI22_X1 U681 ( .A1(n1746), .A2(n6665), .B1(n6042), .B2(n2733), .ZN(n3756)
         );
  OAI22_X1 U682 ( .A1(n1744), .A2(n6666), .B1(n6042), .B2(n2771), .ZN(n3757)
         );
  OAI22_X1 U683 ( .A1(n1742), .A2(n6668), .B1(n6042), .B2(n2734), .ZN(n3758)
         );
  OAI22_X1 U684 ( .A1(n1740), .A2(n6666), .B1(n6042), .B2(n2735), .ZN(n3759)
         );
  OAI22_X1 U685 ( .A1(n1738), .A2(n6671), .B1(n6042), .B2(n2772), .ZN(n3760)
         );
  OAI22_X1 U686 ( .A1(n1736), .A2(n6667), .B1(n6042), .B2(n2736), .ZN(n3761)
         );
  OAI22_X1 U687 ( .A1(n1734), .A2(n6668), .B1(n6042), .B2(n2737), .ZN(n3762)
         );
  OAI22_X1 U688 ( .A1(n1732), .A2(n6668), .B1(n6042), .B2(n2773), .ZN(n3763)
         );
  OAI22_X1 U689 ( .A1(n1730), .A2(n6670), .B1(n6042), .B2(n2738), .ZN(n3764)
         );
  OAI22_X1 U690 ( .A1(n1728), .A2(n6670), .B1(n6042), .B2(n2739), .ZN(n3765)
         );
  OAI22_X1 U691 ( .A1(n1726), .A2(n6669), .B1(n6042), .B2(n2774), .ZN(n3766)
         );
  OAI22_X1 U692 ( .A1(n1724), .A2(n6667), .B1(n6043), .B2(n2740), .ZN(n3767)
         );
  OAI22_X1 U693 ( .A1(n1722), .A2(n6668), .B1(n6043), .B2(n2741), .ZN(n3768)
         );
  OAI22_X1 U694 ( .A1(n1720), .A2(n6667), .B1(n6043), .B2(n2775), .ZN(n3769)
         );
  OAI22_X1 U695 ( .A1(n1718), .A2(n6669), .B1(n6043), .B2(n2742), .ZN(n3770)
         );
  OAI22_X1 U696 ( .A1(n1716), .A2(n6669), .B1(n6043), .B2(n2743), .ZN(n3771)
         );
  OAI22_X1 U697 ( .A1(n1714), .A2(n6669), .B1(n6043), .B2(n2776), .ZN(n3772)
         );
  OAI22_X1 U698 ( .A1(n1712), .A2(n6670), .B1(n6043), .B2(n2744), .ZN(n3773)
         );
  OAI22_X1 U699 ( .A1(n1710), .A2(n6666), .B1(n6043), .B2(n2745), .ZN(n3774)
         );
  OAI22_X1 U700 ( .A1(n1708), .A2(n6670), .B1(n6043), .B2(n2777), .ZN(n3775)
         );
  OAI22_X1 U701 ( .A1(n1706), .A2(n6669), .B1(n6043), .B2(n2746), .ZN(n3776)
         );
  OAI22_X1 U702 ( .A1(n1704), .A2(n6670), .B1(n6043), .B2(n2747), .ZN(n3777)
         );
  OAI22_X1 U703 ( .A1(n1702), .A2(n6671), .B1(n6043), .B2(n2778), .ZN(n3778)
         );
  OAI22_X1 U704 ( .A1(n1748), .A2(n6676), .B1(n6045), .B2(n4325), .ZN(n3787)
         );
  OAI22_X1 U705 ( .A1(n1746), .A2(n6674), .B1(n6045), .B2(n4326), .ZN(n3788)
         );
  OAI22_X1 U706 ( .A1(n1744), .A2(n6676), .B1(n6045), .B2(n5764), .ZN(n3789)
         );
  OAI22_X1 U707 ( .A1(n1742), .A2(n6675), .B1(n6045), .B2(n4327), .ZN(n3790)
         );
  OAI22_X1 U708 ( .A1(n1740), .A2(n6674), .B1(n6045), .B2(n4328), .ZN(n3791)
         );
  OAI22_X1 U709 ( .A1(n1738), .A2(n6679), .B1(n6045), .B2(n5765), .ZN(n3792)
         );
  OAI22_X1 U710 ( .A1(n1736), .A2(n6675), .B1(n6045), .B2(n4329), .ZN(n3793)
         );
  OAI22_X1 U711 ( .A1(n1734), .A2(n6676), .B1(n6045), .B2(n4330), .ZN(n3794)
         );
  OAI22_X1 U712 ( .A1(n1732), .A2(n6676), .B1(n6045), .B2(n5766), .ZN(n3795)
         );
  OAI22_X1 U713 ( .A1(n1730), .A2(n6679), .B1(n6045), .B2(n4331), .ZN(n3796)
         );
  OAI22_X1 U714 ( .A1(n1728), .A2(n6677), .B1(n6045), .B2(n4332), .ZN(n3797)
         );
  OAI22_X1 U715 ( .A1(n1726), .A2(n6678), .B1(n6045), .B2(n5767), .ZN(n3798)
         );
  OAI22_X1 U716 ( .A1(n1724), .A2(n6675), .B1(n6046), .B2(n4333), .ZN(n3799)
         );
  OAI22_X1 U717 ( .A1(n1722), .A2(n6676), .B1(n6046), .B2(n4334), .ZN(n3800)
         );
  OAI22_X1 U718 ( .A1(n1720), .A2(n6675), .B1(n6046), .B2(n5768), .ZN(n3801)
         );
  OAI22_X1 U719 ( .A1(n1718), .A2(n6680), .B1(n6046), .B2(n4335), .ZN(n3802)
         );
  OAI22_X1 U720 ( .A1(n1716), .A2(n6677), .B1(n6046), .B2(n4336), .ZN(n3803)
         );
  OAI22_X1 U721 ( .A1(n1714), .A2(n6678), .B1(n6046), .B2(n5769), .ZN(n3804)
         );
  OAI22_X1 U722 ( .A1(n1712), .A2(n6678), .B1(n6046), .B2(n4337), .ZN(n3805)
         );
  OAI22_X1 U723 ( .A1(n1710), .A2(n6674), .B1(n6046), .B2(n4338), .ZN(n3806)
         );
  OAI22_X1 U724 ( .A1(n1708), .A2(n6677), .B1(n6046), .B2(n5770), .ZN(n3807)
         );
  OAI22_X1 U725 ( .A1(n1706), .A2(n6680), .B1(n6046), .B2(n4339), .ZN(n3808)
         );
  OAI22_X1 U726 ( .A1(n1704), .A2(n6679), .B1(n6046), .B2(n4340), .ZN(n3809)
         );
  OAI22_X1 U727 ( .A1(n1702), .A2(n6680), .B1(n6046), .B2(n5771), .ZN(n3810)
         );
  OAI22_X1 U728 ( .A1(n1748), .A2(n6684), .B1(n6048), .B2(n2792), .ZN(n3819)
         );
  OAI22_X1 U729 ( .A1(n1746), .A2(n6683), .B1(n6048), .B2(n2794), .ZN(n3820)
         );
  OAI22_X1 U730 ( .A1(n1744), .A2(n6684), .B1(n6048), .B2(n2796), .ZN(n3821)
         );
  OAI22_X1 U731 ( .A1(n1742), .A2(n6686), .B1(n6048), .B2(n2798), .ZN(n3822)
         );
  OAI22_X1 U732 ( .A1(n1740), .A2(n6684), .B1(n6048), .B2(n2800), .ZN(n3823)
         );
  OAI22_X1 U733 ( .A1(n1738), .A2(n6689), .B1(n6048), .B2(n2802), .ZN(n3824)
         );
  OAI22_X1 U734 ( .A1(n1736), .A2(n6685), .B1(n6048), .B2(n2804), .ZN(n3825)
         );
  OAI22_X1 U735 ( .A1(n1734), .A2(n6686), .B1(n6048), .B2(n2806), .ZN(n3826)
         );
  OAI22_X1 U736 ( .A1(n1732), .A2(n6686), .B1(n6048), .B2(n2808), .ZN(n3827)
         );
  OAI22_X1 U737 ( .A1(n1730), .A2(n6688), .B1(n6048), .B2(n2810), .ZN(n3828)
         );
  OAI22_X1 U738 ( .A1(n1728), .A2(n6688), .B1(n6048), .B2(n2812), .ZN(n3829)
         );
  OAI22_X1 U739 ( .A1(n1726), .A2(n6687), .B1(n6048), .B2(n2814), .ZN(n3830)
         );
  OAI22_X1 U740 ( .A1(n1724), .A2(n6685), .B1(n6049), .B2(n2816), .ZN(n3831)
         );
  OAI22_X1 U741 ( .A1(n1722), .A2(n6686), .B1(n6049), .B2(n2818), .ZN(n3832)
         );
  OAI22_X1 U742 ( .A1(n1720), .A2(n6685), .B1(n6049), .B2(n2820), .ZN(n3833)
         );
  OAI22_X1 U743 ( .A1(n1718), .A2(n6687), .B1(n6049), .B2(n2822), .ZN(n3834)
         );
  OAI22_X1 U744 ( .A1(n1716), .A2(n6687), .B1(n6049), .B2(n2826), .ZN(n3835)
         );
  OAI22_X1 U745 ( .A1(n1714), .A2(n6687), .B1(n6049), .B2(n2828), .ZN(n3836)
         );
  OAI22_X1 U746 ( .A1(n1712), .A2(n6688), .B1(n6049), .B2(n2830), .ZN(n3837)
         );
  OAI22_X1 U747 ( .A1(n1710), .A2(n6684), .B1(n6049), .B2(n2832), .ZN(n3838)
         );
  OAI22_X1 U748 ( .A1(n1708), .A2(n6688), .B1(n6049), .B2(n2834), .ZN(n3839)
         );
  OAI22_X1 U749 ( .A1(n1706), .A2(n6687), .B1(n6049), .B2(n2836), .ZN(n3840)
         );
  OAI22_X1 U750 ( .A1(n1704), .A2(n6688), .B1(n6049), .B2(n2838), .ZN(n3841)
         );
  OAI22_X1 U751 ( .A1(n1702), .A2(n6689), .B1(n6049), .B2(n2839), .ZN(n3842)
         );
  OAI22_X1 U752 ( .A1(n1748), .A2(n6694), .B1(n6051), .B2(n5784), .ZN(n3851)
         );
  OAI22_X1 U753 ( .A1(n1746), .A2(n6692), .B1(n6051), .B2(n5786), .ZN(n3852)
         );
  OAI22_X1 U754 ( .A1(n1744), .A2(n6694), .B1(n6051), .B2(n5788), .ZN(n3853)
         );
  OAI22_X1 U755 ( .A1(n1742), .A2(n6693), .B1(n6051), .B2(n5790), .ZN(n3854)
         );
  OAI22_X1 U756 ( .A1(n1740), .A2(n6692), .B1(n6051), .B2(n5792), .ZN(n3855)
         );
  OAI22_X1 U757 ( .A1(n1738), .A2(n6697), .B1(n6051), .B2(n5794), .ZN(n3856)
         );
  OAI22_X1 U758 ( .A1(n1736), .A2(n6693), .B1(n6051), .B2(n5796), .ZN(n3857)
         );
  OAI22_X1 U759 ( .A1(n1734), .A2(n6694), .B1(n6051), .B2(n5798), .ZN(n3858)
         );
  OAI22_X1 U760 ( .A1(n1732), .A2(n6694), .B1(n6051), .B2(n5800), .ZN(n3859)
         );
  OAI22_X1 U761 ( .A1(n1730), .A2(n6697), .B1(n6051), .B2(n5802), .ZN(n3860)
         );
  OAI22_X1 U762 ( .A1(n1728), .A2(n6695), .B1(n6051), .B2(n5804), .ZN(n3861)
         );
  OAI22_X1 U763 ( .A1(n1726), .A2(n6696), .B1(n6051), .B2(n5806), .ZN(n3862)
         );
  OAI22_X1 U764 ( .A1(n1724), .A2(n6693), .B1(n6052), .B2(n5808), .ZN(n3863)
         );
  OAI22_X1 U765 ( .A1(n1722), .A2(n6694), .B1(n6052), .B2(n5810), .ZN(n3864)
         );
  OAI22_X1 U766 ( .A1(n1720), .A2(n6693), .B1(n6052), .B2(n5812), .ZN(n3865)
         );
  OAI22_X1 U767 ( .A1(n1718), .A2(n6698), .B1(n6052), .B2(n5814), .ZN(n3866)
         );
  OAI22_X1 U768 ( .A1(n1716), .A2(n6695), .B1(n6052), .B2(n5816), .ZN(n3867)
         );
  OAI22_X1 U769 ( .A1(n1714), .A2(n6696), .B1(n6052), .B2(n5818), .ZN(n3868)
         );
  OAI22_X1 U770 ( .A1(n1712), .A2(n6696), .B1(n6052), .B2(n5820), .ZN(n3869)
         );
  OAI22_X1 U771 ( .A1(n1710), .A2(n6692), .B1(n6052), .B2(n5822), .ZN(n3870)
         );
  OAI22_X1 U772 ( .A1(n1708), .A2(n6695), .B1(n6052), .B2(n5824), .ZN(n3871)
         );
  OAI22_X1 U773 ( .A1(n1706), .A2(n6698), .B1(n6052), .B2(n5826), .ZN(n3872)
         );
  OAI22_X1 U774 ( .A1(n1704), .A2(n6697), .B1(n6052), .B2(n5828), .ZN(n3873)
         );
  OAI22_X1 U775 ( .A1(n1702), .A2(n6698), .B1(n6052), .B2(n5829), .ZN(n3874)
         );
  OAI22_X1 U776 ( .A1(n1748), .A2(n6732), .B1(n6066), .B2(n4296), .ZN(n4011)
         );
  OAI22_X1 U777 ( .A1(n1746), .A2(n1822), .B1(n6066), .B2(n4297), .ZN(n4012)
         );
  OAI22_X1 U778 ( .A1(n1744), .A2(n6731), .B1(n6066), .B2(n4298), .ZN(n4013)
         );
  OAI22_X1 U779 ( .A1(n1742), .A2(n6732), .B1(n6066), .B2(n4299), .ZN(n4014)
         );
  OAI22_X1 U780 ( .A1(n1740), .A2(n1822), .B1(n6066), .B2(n4300), .ZN(n4015)
         );
  OAI22_X1 U781 ( .A1(n1738), .A2(n6731), .B1(n6066), .B2(n4301), .ZN(n4016)
         );
  OAI22_X1 U782 ( .A1(n1736), .A2(n6732), .B1(n6066), .B2(n4302), .ZN(n4017)
         );
  OAI22_X1 U783 ( .A1(n1734), .A2(n1822), .B1(n6066), .B2(n4303), .ZN(n4018)
         );
  OAI22_X1 U784 ( .A1(n1732), .A2(n6731), .B1(n6066), .B2(n4304), .ZN(n4019)
         );
  OAI22_X1 U785 ( .A1(n1730), .A2(n6732), .B1(n6066), .B2(n4305), .ZN(n4020)
         );
  OAI22_X1 U786 ( .A1(n1728), .A2(n1822), .B1(n6066), .B2(n4306), .ZN(n4021)
         );
  OAI22_X1 U787 ( .A1(n1726), .A2(n6731), .B1(n6066), .B2(n4307), .ZN(n4022)
         );
  OAI22_X1 U788 ( .A1(n1724), .A2(n6732), .B1(n6067), .B2(n4308), .ZN(n4023)
         );
  OAI22_X1 U789 ( .A1(n1722), .A2(n1822), .B1(n6067), .B2(n4309), .ZN(n4024)
         );
  OAI22_X1 U790 ( .A1(n1720), .A2(n6731), .B1(n6067), .B2(n4310), .ZN(n4025)
         );
  OAI22_X1 U791 ( .A1(n1718), .A2(n6732), .B1(n6067), .B2(n4311), .ZN(n4026)
         );
  OAI22_X1 U792 ( .A1(n1716), .A2(n1822), .B1(n6067), .B2(n4312), .ZN(n4027)
         );
  OAI22_X1 U793 ( .A1(n1714), .A2(n6731), .B1(n6067), .B2(n4313), .ZN(n4028)
         );
  OAI22_X1 U794 ( .A1(n1712), .A2(n6732), .B1(n6067), .B2(n4314), .ZN(n4029)
         );
  OAI22_X1 U795 ( .A1(n1710), .A2(n1822), .B1(n6067), .B2(n4315), .ZN(n4030)
         );
  OAI22_X1 U796 ( .A1(n1708), .A2(n6731), .B1(n6067), .B2(n4316), .ZN(n4031)
         );
  OAI22_X1 U797 ( .A1(n1706), .A2(n6732), .B1(n6067), .B2(n4317), .ZN(n4032)
         );
  OAI22_X1 U798 ( .A1(n1704), .A2(n1822), .B1(n6067), .B2(n5901), .ZN(n4033)
         );
  OAI22_X1 U799 ( .A1(n1702), .A2(n6731), .B1(n6067), .B2(n5903), .ZN(n4034)
         );
  OAI22_X1 U800 ( .A1(n1748), .A2(n6734), .B1(n6069), .B2(n2569), .ZN(n4043)
         );
  OAI22_X1 U801 ( .A1(n1746), .A2(n1787), .B1(n6069), .B2(n2570), .ZN(n4044)
         );
  OAI22_X1 U802 ( .A1(n1744), .A2(n6733), .B1(n6069), .B2(n2571), .ZN(n4045)
         );
  OAI22_X1 U803 ( .A1(n1742), .A2(n6734), .B1(n6069), .B2(n2572), .ZN(n4046)
         );
  OAI22_X1 U804 ( .A1(n1740), .A2(n1787), .B1(n6069), .B2(n2573), .ZN(n4047)
         );
  OAI22_X1 U805 ( .A1(n1738), .A2(n6733), .B1(n6069), .B2(n2574), .ZN(n4048)
         );
  OAI22_X1 U806 ( .A1(n1736), .A2(n6734), .B1(n6069), .B2(n2575), .ZN(n4049)
         );
  OAI22_X1 U807 ( .A1(n1734), .A2(n1787), .B1(n6069), .B2(n2576), .ZN(n4050)
         );
  OAI22_X1 U808 ( .A1(n1732), .A2(n6733), .B1(n6069), .B2(n2577), .ZN(n4051)
         );
  OAI22_X1 U809 ( .A1(n1730), .A2(n6734), .B1(n6069), .B2(n2578), .ZN(n4052)
         );
  OAI22_X1 U810 ( .A1(n1728), .A2(n1787), .B1(n6069), .B2(n2579), .ZN(n4053)
         );
  OAI22_X1 U811 ( .A1(n1726), .A2(n6733), .B1(n6069), .B2(n2580), .ZN(n4054)
         );
  OAI22_X1 U812 ( .A1(n1724), .A2(n6734), .B1(n6070), .B2(n2581), .ZN(n4055)
         );
  OAI22_X1 U813 ( .A1(n1722), .A2(n1787), .B1(n6070), .B2(n2583), .ZN(n4056)
         );
  OAI22_X1 U814 ( .A1(n1720), .A2(n6733), .B1(n6070), .B2(n2618), .ZN(n4057)
         );
  OAI22_X1 U815 ( .A1(n1718), .A2(n6734), .B1(n6070), .B2(n2652), .ZN(n4058)
         );
  OAI22_X1 U816 ( .A1(n1716), .A2(n1787), .B1(n6070), .B2(n2686), .ZN(n4059)
         );
  OAI22_X1 U817 ( .A1(n1714), .A2(n6733), .B1(n6070), .B2(n2723), .ZN(n4060)
         );
  OAI22_X1 U818 ( .A1(n1712), .A2(n6734), .B1(n6070), .B2(n2724), .ZN(n4061)
         );
  OAI22_X1 U819 ( .A1(n1710), .A2(n1787), .B1(n6070), .B2(n2725), .ZN(n4062)
         );
  OAI22_X1 U820 ( .A1(n1708), .A2(n6733), .B1(n6070), .B2(n2726), .ZN(n4063)
         );
  OAI22_X1 U821 ( .A1(n1706), .A2(n6734), .B1(n6070), .B2(n2727), .ZN(n4064)
         );
  OAI22_X1 U822 ( .A1(n1704), .A2(n1787), .B1(n6070), .B2(n4202), .ZN(n4065)
         );
  OAI22_X1 U823 ( .A1(n1702), .A2(n6733), .B1(n6070), .B2(n4204), .ZN(n4066)
         );
  NAND2_X1 U824 ( .A1(n5732), .A2(n5724), .ZN(n5115) );
  NAND2_X1 U825 ( .A1(n5733), .A2(n5724), .ZN(n5114) );
  OAI22_X1 U826 ( .A1(n1700), .A2(n6513), .B1(n5990), .B2(n4272), .ZN(n3203)
         );
  OAI22_X1 U827 ( .A1(n1698), .A2(n6514), .B1(n5990), .B2(n4273), .ZN(n3204)
         );
  OAI22_X1 U828 ( .A1(n1696), .A2(n6516), .B1(n5990), .B2(n4274), .ZN(n3205)
         );
  OAI22_X1 U829 ( .A1(n1694), .A2(n6516), .B1(n5990), .B2(n4275), .ZN(n3206)
         );
  OAI22_X1 U830 ( .A1(n1692), .A2(n6516), .B1(n5990), .B2(n4276), .ZN(n3207)
         );
  OAI22_X1 U831 ( .A1(n1690), .A2(n6516), .B1(n5990), .B2(n4277), .ZN(n3208)
         );
  OAI22_X1 U832 ( .A1(n1688), .A2(n6511), .B1(n5990), .B2(n4278), .ZN(n3209)
         );
  OAI22_X1 U833 ( .A1(n1685), .A2(n6515), .B1(n5990), .B2(n4279), .ZN(n3210)
         );
  OAI22_X1 U834 ( .A1(n1700), .A2(n6524), .B1(n5993), .B2(n5968), .ZN(n3235)
         );
  OAI22_X1 U835 ( .A1(n1698), .A2(n6520), .B1(n5993), .B2(n5969), .ZN(n3236)
         );
  OAI22_X1 U836 ( .A1(n1696), .A2(n6521), .B1(n5993), .B2(n5970), .ZN(n3237)
         );
  OAI22_X1 U837 ( .A1(n1694), .A2(n6521), .B1(n5993), .B2(n5971), .ZN(n3238)
         );
  OAI22_X1 U838 ( .A1(n1692), .A2(n6522), .B1(n5993), .B2(n5972), .ZN(n3239)
         );
  OAI22_X1 U839 ( .A1(n1690), .A2(n6523), .B1(n5993), .B2(n5973), .ZN(n3240)
         );
  OAI22_X1 U840 ( .A1(n1688), .A2(n6524), .B1(n5993), .B2(n5974), .ZN(n3241)
         );
  OAI22_X1 U841 ( .A1(n1685), .A2(n6524), .B1(n5993), .B2(n5975), .ZN(n3242)
         );
  OAI22_X1 U842 ( .A1(n1700), .A2(n6529), .B1(n5996), .B2(n4205), .ZN(n3267)
         );
  OAI22_X1 U843 ( .A1(n1698), .A2(n6530), .B1(n5996), .B2(n4207), .ZN(n3268)
         );
  OAI22_X1 U844 ( .A1(n1696), .A2(n6532), .B1(n5996), .B2(n4209), .ZN(n3269)
         );
  OAI22_X1 U845 ( .A1(n1694), .A2(n6532), .B1(n5996), .B2(n4211), .ZN(n3270)
         );
  OAI22_X1 U846 ( .A1(n1692), .A2(n6532), .B1(n5996), .B2(n4191), .ZN(n3271)
         );
  OAI22_X1 U847 ( .A1(n1690), .A2(n6532), .B1(n5996), .B2(n4193), .ZN(n3272)
         );
  OAI22_X1 U848 ( .A1(n1688), .A2(n6527), .B1(n5996), .B2(n4195), .ZN(n3273)
         );
  OAI22_X1 U849 ( .A1(n1685), .A2(n6531), .B1(n5996), .B2(n4197), .ZN(n3274)
         );
  OAI22_X1 U850 ( .A1(n1700), .A2(n6541), .B1(n5999), .B2(n5904), .ZN(n3299)
         );
  OAI22_X1 U851 ( .A1(n1698), .A2(n6541), .B1(n5999), .B2(n5906), .ZN(n3300)
         );
  OAI22_X1 U852 ( .A1(n1696), .A2(n6537), .B1(n5999), .B2(n5908), .ZN(n3301)
         );
  OAI22_X1 U853 ( .A1(n1694), .A2(n6538), .B1(n5999), .B2(n5910), .ZN(n3302)
         );
  OAI22_X1 U854 ( .A1(n1692), .A2(n6534), .B1(n5999), .B2(n5890), .ZN(n3303)
         );
  OAI22_X1 U855 ( .A1(n1690), .A2(n6535), .B1(n5999), .B2(n5892), .ZN(n3304)
         );
  OAI22_X1 U856 ( .A1(n1688), .A2(n6537), .B1(n5999), .B2(n5894), .ZN(n3305)
         );
  OAI22_X1 U857 ( .A1(n1685), .A2(n6536), .B1(n5999), .B2(n5896), .ZN(n3306)
         );
  OAI22_X1 U858 ( .A1(n1700), .A2(n6546), .B1(n6002), .B2(n4282), .ZN(n3331)
         );
  OAI22_X1 U859 ( .A1(n1698), .A2(n6547), .B1(n6002), .B2(n4283), .ZN(n3332)
         );
  OAI22_X1 U860 ( .A1(n1696), .A2(n6549), .B1(n6002), .B2(n4284), .ZN(n3333)
         );
  OAI22_X1 U861 ( .A1(n1694), .A2(n6549), .B1(n6002), .B2(n4287), .ZN(n3334)
         );
  OAI22_X1 U862 ( .A1(n1692), .A2(n6549), .B1(n6002), .B2(n4242), .ZN(n3335)
         );
  OAI22_X1 U863 ( .A1(n1690), .A2(n6549), .B1(n6002), .B2(n4243), .ZN(n3336)
         );
  OAI22_X1 U864 ( .A1(n1688), .A2(n6544), .B1(n6002), .B2(n4244), .ZN(n3337)
         );
  OAI22_X1 U865 ( .A1(n1685), .A2(n6548), .B1(n6002), .B2(n4245), .ZN(n3338)
         );
  OAI22_X1 U866 ( .A1(n1700), .A2(n6557), .B1(n6005), .B2(n5978), .ZN(n3363)
         );
  OAI22_X1 U867 ( .A1(n1698), .A2(n6553), .B1(n6005), .B2(n5979), .ZN(n3364)
         );
  OAI22_X1 U868 ( .A1(n1696), .A2(n6554), .B1(n6005), .B2(n5980), .ZN(n3365)
         );
  OAI22_X1 U869 ( .A1(n1694), .A2(n6554), .B1(n6005), .B2(n5981), .ZN(n3366)
         );
  OAI22_X1 U870 ( .A1(n1692), .A2(n6555), .B1(n6005), .B2(n5940), .ZN(n3367)
         );
  OAI22_X1 U871 ( .A1(n1690), .A2(n6556), .B1(n6005), .B2(n5941), .ZN(n3368)
         );
  OAI22_X1 U872 ( .A1(n1688), .A2(n6557), .B1(n6005), .B2(n5942), .ZN(n3369)
         );
  OAI22_X1 U873 ( .A1(n1685), .A2(n6557), .B1(n6005), .B2(n5943), .ZN(n3370)
         );
  OAI22_X1 U874 ( .A1(n1700), .A2(n6598), .B1(n6020), .B2(n4187), .ZN(n3523)
         );
  OAI22_X1 U875 ( .A1(n1698), .A2(n6599), .B1(n6020), .B2(n4188), .ZN(n3524)
         );
  OAI22_X1 U876 ( .A1(n1696), .A2(n6601), .B1(n6020), .B2(n4189), .ZN(n3525)
         );
  OAI22_X1 U877 ( .A1(n1694), .A2(n6601), .B1(n6020), .B2(n4190), .ZN(n3526)
         );
  OAI22_X1 U878 ( .A1(n1692), .A2(n6601), .B1(n6020), .B2(n4192), .ZN(n3527)
         );
  OAI22_X1 U879 ( .A1(n1690), .A2(n6601), .B1(n6020), .B2(n4194), .ZN(n3528)
         );
  OAI22_X1 U880 ( .A1(n1688), .A2(n6596), .B1(n6020), .B2(n4196), .ZN(n3529)
         );
  OAI22_X1 U881 ( .A1(n1685), .A2(n6600), .B1(n6020), .B2(n4198), .ZN(n3530)
         );
  OAI22_X1 U882 ( .A1(n1700), .A2(n6610), .B1(n6023), .B2(n5886), .ZN(n3555)
         );
  OAI22_X1 U883 ( .A1(n1698), .A2(n6610), .B1(n6023), .B2(n5887), .ZN(n3556)
         );
  OAI22_X1 U884 ( .A1(n1696), .A2(n6606), .B1(n6023), .B2(n5888), .ZN(n3557)
         );
  OAI22_X1 U885 ( .A1(n1694), .A2(n6607), .B1(n6023), .B2(n5889), .ZN(n3558)
         );
  OAI22_X1 U886 ( .A1(n1692), .A2(n6603), .B1(n6023), .B2(n5891), .ZN(n3559)
         );
  OAI22_X1 U887 ( .A1(n1690), .A2(n6604), .B1(n6023), .B2(n5893), .ZN(n3560)
         );
  OAI22_X1 U888 ( .A1(n1688), .A2(n6606), .B1(n6023), .B2(n5895), .ZN(n3561)
         );
  OAI22_X1 U889 ( .A1(n1685), .A2(n6605), .B1(n6023), .B2(n5897), .ZN(n3562)
         );
  OAI22_X1 U890 ( .A1(n1700), .A2(n6615), .B1(n6026), .B2(n4215), .ZN(n3587)
         );
  OAI22_X1 U891 ( .A1(n1698), .A2(n6616), .B1(n6026), .B2(n4216), .ZN(n3588)
         );
  OAI22_X1 U892 ( .A1(n1696), .A2(n6618), .B1(n6026), .B2(n4218), .ZN(n3589)
         );
  OAI22_X1 U893 ( .A1(n1694), .A2(n6618), .B1(n6026), .B2(n4219), .ZN(n3590)
         );
  OAI22_X1 U894 ( .A1(n1692), .A2(n6618), .B1(n6026), .B2(n2845), .ZN(n3591)
         );
  OAI22_X1 U895 ( .A1(n1690), .A2(n6618), .B1(n6026), .B2(n2847), .ZN(n3592)
         );
  OAI22_X1 U896 ( .A1(n1688), .A2(n6613), .B1(n6026), .B2(n2849), .ZN(n3593)
         );
  OAI22_X1 U897 ( .A1(n1685), .A2(n6617), .B1(n6026), .B2(n2851), .ZN(n3594)
         );
  OAI22_X1 U898 ( .A1(n1700), .A2(n6626), .B1(n6029), .B2(n5914), .ZN(n3619)
         );
  OAI22_X1 U899 ( .A1(n1698), .A2(n6622), .B1(n6029), .B2(n5915), .ZN(n3620)
         );
  OAI22_X1 U900 ( .A1(n1696), .A2(n6623), .B1(n6029), .B2(n5916), .ZN(n3621)
         );
  OAI22_X1 U901 ( .A1(n1694), .A2(n6623), .B1(n6029), .B2(n5917), .ZN(n3622)
         );
  OAI22_X1 U902 ( .A1(n1692), .A2(n6624), .B1(n6029), .B2(n5835), .ZN(n3623)
         );
  OAI22_X1 U903 ( .A1(n1690), .A2(n6625), .B1(n6029), .B2(n5837), .ZN(n3624)
         );
  OAI22_X1 U904 ( .A1(n1688), .A2(n6626), .B1(n6029), .B2(n5839), .ZN(n3625)
         );
  OAI22_X1 U905 ( .A1(n1685), .A2(n6626), .B1(n6029), .B2(n5841), .ZN(n3626)
         );
  OAI22_X1 U906 ( .A1(n1700), .A2(n6671), .B1(n6044), .B2(n2748), .ZN(n3779)
         );
  OAI22_X1 U907 ( .A1(n1698), .A2(n6671), .B1(n6044), .B2(n2749), .ZN(n3780)
         );
  OAI22_X1 U908 ( .A1(n1696), .A2(n6671), .B1(n6044), .B2(n2779), .ZN(n3781)
         );
  OAI22_X1 U909 ( .A1(n1694), .A2(n6671), .B1(n6044), .B2(n2750), .ZN(n3782)
         );
  OAI22_X1 U910 ( .A1(n1692), .A2(n6665), .B1(n6044), .B2(n2751), .ZN(n3783)
         );
  OAI22_X1 U911 ( .A1(n1690), .A2(n6665), .B1(n6044), .B2(n2780), .ZN(n3784)
         );
  OAI22_X1 U912 ( .A1(n1688), .A2(n6665), .B1(n6044), .B2(n2752), .ZN(n3785)
         );
  OAI22_X1 U913 ( .A1(n1685), .A2(n6667), .B1(n6044), .B2(n2753), .ZN(n3786)
         );
  OAI22_X1 U914 ( .A1(n1700), .A2(n6679), .B1(n6047), .B2(n4341), .ZN(n3811)
         );
  OAI22_X1 U915 ( .A1(n1698), .A2(n6679), .B1(n6047), .B2(n4342), .ZN(n3812)
         );
  OAI22_X1 U916 ( .A1(n1696), .A2(n6680), .B1(n6047), .B2(n5772), .ZN(n3813)
         );
  OAI22_X1 U917 ( .A1(n1694), .A2(n6680), .B1(n6047), .B2(n4343), .ZN(n3814)
         );
  OAI22_X1 U918 ( .A1(n1692), .A2(n6676), .B1(n6047), .B2(n4344), .ZN(n3815)
         );
  OAI22_X1 U919 ( .A1(n1690), .A2(n6675), .B1(n6047), .B2(n5773), .ZN(n3816)
         );
  OAI22_X1 U920 ( .A1(n1688), .A2(n6678), .B1(n6047), .B2(n4345), .ZN(n3817)
         );
  OAI22_X1 U921 ( .A1(n1685), .A2(n6677), .B1(n6047), .B2(n4346), .ZN(n3818)
         );
  OAI22_X1 U922 ( .A1(n1700), .A2(n6689), .B1(n6050), .B2(n2840), .ZN(n3843)
         );
  OAI22_X1 U923 ( .A1(n1698), .A2(n6689), .B1(n6050), .B2(n2841), .ZN(n3844)
         );
  OAI22_X1 U924 ( .A1(n1696), .A2(n6689), .B1(n6050), .B2(n2842), .ZN(n3845)
         );
  OAI22_X1 U925 ( .A1(n1694), .A2(n6689), .B1(n6050), .B2(n2843), .ZN(n3846)
         );
  OAI22_X1 U926 ( .A1(n1692), .A2(n6683), .B1(n6050), .B2(n2844), .ZN(n3847)
         );
  OAI22_X1 U927 ( .A1(n1690), .A2(n6683), .B1(n6050), .B2(n2846), .ZN(n3848)
         );
  OAI22_X1 U928 ( .A1(n1688), .A2(n6683), .B1(n6050), .B2(n2848), .ZN(n3849)
         );
  OAI22_X1 U929 ( .A1(n1685), .A2(n6685), .B1(n6050), .B2(n2850), .ZN(n3850)
         );
  OAI22_X1 U930 ( .A1(n1700), .A2(n6697), .B1(n6053), .B2(n5830), .ZN(n3875)
         );
  OAI22_X1 U931 ( .A1(n1698), .A2(n6697), .B1(n6053), .B2(n5831), .ZN(n3876)
         );
  OAI22_X1 U932 ( .A1(n1696), .A2(n6698), .B1(n6053), .B2(n5832), .ZN(n3877)
         );
  OAI22_X1 U933 ( .A1(n1694), .A2(n6698), .B1(n6053), .B2(n5833), .ZN(n3878)
         );
  OAI22_X1 U934 ( .A1(n1692), .A2(n6694), .B1(n6053), .B2(n5834), .ZN(n3879)
         );
  OAI22_X1 U935 ( .A1(n1690), .A2(n6693), .B1(n6053), .B2(n5836), .ZN(n3880)
         );
  OAI22_X1 U936 ( .A1(n1688), .A2(n6696), .B1(n6053), .B2(n5838), .ZN(n3881)
         );
  OAI22_X1 U937 ( .A1(n1685), .A2(n6695), .B1(n6053), .B2(n5840), .ZN(n3882)
         );
  OAI22_X1 U938 ( .A1(n1700), .A2(n6732), .B1(n6068), .B2(n5905), .ZN(n4035)
         );
  OAI22_X1 U939 ( .A1(n1698), .A2(n1822), .B1(n6068), .B2(n5907), .ZN(n4036)
         );
  OAI22_X1 U940 ( .A1(n1696), .A2(n6731), .B1(n6068), .B2(n5909), .ZN(n4037)
         );
  OAI22_X1 U941 ( .A1(n1694), .A2(n6732), .B1(n6068), .B2(n5911), .ZN(n4038)
         );
  OAI22_X1 U942 ( .A1(n1692), .A2(n1822), .B1(n6068), .B2(n4318), .ZN(n4039)
         );
  OAI22_X1 U943 ( .A1(n1690), .A2(n6731), .B1(n6068), .B2(n4322), .ZN(n4040)
         );
  OAI22_X1 U944 ( .A1(n1688), .A2(n6732), .B1(n6068), .B2(n4323), .ZN(n4041)
         );
  OAI22_X1 U945 ( .A1(n1685), .A2(n1822), .B1(n6068), .B2(n4324), .ZN(n4042)
         );
  OAI22_X1 U946 ( .A1(n1700), .A2(n6734), .B1(n6071), .B2(n4206), .ZN(n4067)
         );
  OAI22_X1 U947 ( .A1(n1698), .A2(n1787), .B1(n6071), .B2(n4208), .ZN(n4068)
         );
  OAI22_X1 U948 ( .A1(n1696), .A2(n6733), .B1(n6071), .B2(n4210), .ZN(n4069)
         );
  OAI22_X1 U949 ( .A1(n1694), .A2(n6734), .B1(n6071), .B2(n4212), .ZN(n4070)
         );
  OAI22_X1 U950 ( .A1(n1692), .A2(n1787), .B1(n6071), .B2(n2728), .ZN(n4071)
         );
  OAI22_X1 U951 ( .A1(n1690), .A2(n6733), .B1(n6071), .B2(n2729), .ZN(n4072)
         );
  OAI22_X1 U952 ( .A1(n1688), .A2(n6734), .B1(n6071), .B2(n2730), .ZN(n4073)
         );
  OAI22_X1 U953 ( .A1(n1685), .A2(n1787), .B1(n6071), .B2(n2731), .ZN(n4074)
         );
  OAI22_X1 U954 ( .A1(n1748), .A2(n6735), .B1(n6744), .B2(n2561), .ZN(n4075)
         );
  OAI22_X1 U955 ( .A1(n1746), .A2(n6735), .B1(n6744), .B2(n2562), .ZN(n4076)
         );
  OAI22_X1 U956 ( .A1(n1744), .A2(n6735), .B1(n6744), .B2(n2781), .ZN(n4077)
         );
  OAI22_X1 U957 ( .A1(n1742), .A2(n6735), .B1(n6744), .B2(n2563), .ZN(n4078)
         );
  OAI22_X1 U958 ( .A1(n1740), .A2(n6735), .B1(n6743), .B2(n2754), .ZN(n4079)
         );
  OAI22_X1 U959 ( .A1(n1738), .A2(n6735), .B1(n6743), .B2(n2782), .ZN(n4080)
         );
  OAI22_X1 U960 ( .A1(n1736), .A2(n6735), .B1(n6743), .B2(n2758), .ZN(n4081)
         );
  OAI22_X1 U961 ( .A1(n1734), .A2(n6735), .B1(n6743), .B2(n2759), .ZN(n4082)
         );
  OAI22_X1 U962 ( .A1(n1732), .A2(n6735), .B1(n6742), .B2(n2783), .ZN(n4083)
         );
  OAI22_X1 U963 ( .A1(n1730), .A2(n6735), .B1(n6742), .B2(n2760), .ZN(n4084)
         );
  OAI22_X1 U964 ( .A1(n1728), .A2(n6735), .B1(n6742), .B2(n2564), .ZN(n4085)
         );
  OAI22_X1 U965 ( .A1(n1726), .A2(n6735), .B1(n6742), .B2(n2784), .ZN(n4086)
         );
  OAI22_X1 U966 ( .A1(n1724), .A2(n6736), .B1(n6741), .B2(n2761), .ZN(n4087)
         );
  OAI22_X1 U967 ( .A1(n1722), .A2(n6736), .B1(n6741), .B2(n2762), .ZN(n4088)
         );
  OAI22_X1 U968 ( .A1(n1720), .A2(n6736), .B1(n6741), .B2(n2785), .ZN(n4089)
         );
  OAI22_X1 U969 ( .A1(n1718), .A2(n6736), .B1(n6741), .B2(n2763), .ZN(n4090)
         );
  OAI22_X1 U970 ( .A1(n1716), .A2(n6736), .B1(n6740), .B2(n2764), .ZN(n4091)
         );
  OAI22_X1 U971 ( .A1(n1714), .A2(n6736), .B1(n6740), .B2(n2786), .ZN(n4092)
         );
  OAI22_X1 U972 ( .A1(n1712), .A2(n6736), .B1(n6740), .B2(n2565), .ZN(n4093)
         );
  OAI22_X1 U973 ( .A1(n1710), .A2(n6736), .B1(n6740), .B2(n2566), .ZN(n4094)
         );
  OAI22_X1 U974 ( .A1(n1708), .A2(n6736), .B1(n6739), .B2(n2787), .ZN(n4095)
         );
  OAI22_X1 U975 ( .A1(n1706), .A2(n6736), .B1(n6739), .B2(n2567), .ZN(n4096)
         );
  OAI22_X1 U976 ( .A1(n1704), .A2(n6736), .B1(n6739), .B2(n2765), .ZN(n4097)
         );
  OAI22_X1 U977 ( .A1(n1702), .A2(n6736), .B1(n6739), .B2(n2788), .ZN(n4098)
         );
  OAI22_X1 U978 ( .A1(n1700), .A2(n6735), .B1(n6738), .B2(n2766), .ZN(n4099)
         );
  OAI22_X1 U979 ( .A1(n1698), .A2(n6736), .B1(n6738), .B2(n2767), .ZN(n4100)
         );
  OAI22_X1 U980 ( .A1(n1696), .A2(n6735), .B1(n6738), .B2(n2789), .ZN(n4101)
         );
  OAI22_X1 U981 ( .A1(n1694), .A2(n6736), .B1(n6738), .B2(n2768), .ZN(n4102)
         );
  OAI22_X1 U982 ( .A1(n1692), .A2(n6735), .B1(n6737), .B2(n2568), .ZN(n4103)
         );
  OAI22_X1 U983 ( .A1(n1690), .A2(n6736), .B1(n6737), .B2(n2791), .ZN(n4104)
         );
  OAI22_X1 U984 ( .A1(n1688), .A2(n6735), .B1(n6737), .B2(n2769), .ZN(n4105)
         );
  OAI22_X1 U985 ( .A1(n1685), .A2(n6736), .B1(n6737), .B2(n2770), .ZN(n4106)
         );
  OAI22_X1 U986 ( .A1(n6749), .A2(n1700), .B1(n6746), .B2(n5759), .ZN(n4131)
         );
  OAI22_X1 U987 ( .A1(n6749), .A2(n1698), .B1(n6747), .B2(n5760), .ZN(n4132)
         );
  OAI22_X1 U988 ( .A1(n6749), .A2(n1696), .B1(n6746), .B2(n5782), .ZN(n4133)
         );
  OAI22_X1 U989 ( .A1(n6748), .A2(n1694), .B1(n6747), .B2(n5761), .ZN(n4134)
         );
  OAI22_X1 U990 ( .A1(n6748), .A2(n1692), .B1(n6746), .B2(n4295), .ZN(n4135)
         );
  OAI22_X1 U991 ( .A1(n6748), .A2(n1690), .B1(n6747), .B2(n5783), .ZN(n4136)
         );
  OAI22_X1 U992 ( .A1(n6748), .A2(n1688), .B1(n6746), .B2(n5762), .ZN(n4137)
         );
  OAI22_X1 U993 ( .A1(n6748), .A2(n1685), .B1(n6747), .B2(n5763), .ZN(n4138)
         );
  OAI22_X1 U994 ( .A1(n6754), .A2(n1748), .B1(n6746), .B2(n4288), .ZN(n4107)
         );
  OAI22_X1 U995 ( .A1(n6754), .A2(n1746), .B1(n6746), .B2(n4289), .ZN(n4108)
         );
  OAI22_X1 U996 ( .A1(n6753), .A2(n1744), .B1(n6746), .B2(n5774), .ZN(n4109)
         );
  OAI22_X1 U997 ( .A1(n6753), .A2(n1742), .B1(n6746), .B2(n4290), .ZN(n4110)
         );
  OAI22_X1 U998 ( .A1(n6753), .A2(n1740), .B1(n6746), .B2(n4347), .ZN(n4111)
         );
  OAI22_X1 U999 ( .A1(n6753), .A2(n1738), .B1(n6746), .B2(n5775), .ZN(n4112)
         );
  OAI22_X1 U1000 ( .A1(n6753), .A2(n1736), .B1(n6746), .B2(n4348), .ZN(n4113)
         );
  OAI22_X1 U1001 ( .A1(n6752), .A2(n1734), .B1(n6746), .B2(n4349), .ZN(n4114)
         );
  OAI22_X1 U1002 ( .A1(n6752), .A2(n1732), .B1(n6746), .B2(n5776), .ZN(n4115)
         );
  OAI22_X1 U1003 ( .A1(n6752), .A2(n1730), .B1(n6746), .B2(n4350), .ZN(n4116)
         );
  OAI22_X1 U1004 ( .A1(n6752), .A2(n1728), .B1(n6746), .B2(n4291), .ZN(n4117)
         );
  OAI22_X1 U1005 ( .A1(n6752), .A2(n1726), .B1(n6746), .B2(n5777), .ZN(n4118)
         );
  OAI22_X1 U1006 ( .A1(n6751), .A2(n1724), .B1(n6747), .B2(n4351), .ZN(n4119)
         );
  OAI22_X1 U1007 ( .A1(n6751), .A2(n1722), .B1(n6747), .B2(n4352), .ZN(n4120)
         );
  OAI22_X1 U1008 ( .A1(n6751), .A2(n1720), .B1(n6747), .B2(n5778), .ZN(n4121)
         );
  OAI22_X1 U1009 ( .A1(n6751), .A2(n1718), .B1(n6747), .B2(n4353), .ZN(n4122)
         );
  OAI22_X1 U1010 ( .A1(n6751), .A2(n1716), .B1(n6747), .B2(n4356), .ZN(n4123)
         );
  OAI22_X1 U1011 ( .A1(n6750), .A2(n1714), .B1(n6747), .B2(n5779), .ZN(n4124)
         );
  OAI22_X1 U1012 ( .A1(n6750), .A2(n1712), .B1(n6747), .B2(n4292), .ZN(n4125)
         );
  OAI22_X1 U1013 ( .A1(n6750), .A2(n1710), .B1(n6747), .B2(n4293), .ZN(n4126)
         );
  OAI22_X1 U1014 ( .A1(n6750), .A2(n1708), .B1(n6747), .B2(n5780), .ZN(n4127)
         );
  OAI22_X1 U1015 ( .A1(n6750), .A2(n1706), .B1(n6747), .B2(n4294), .ZN(n4128)
         );
  OAI22_X1 U1016 ( .A1(n6749), .A2(n1704), .B1(n6747), .B2(n4390), .ZN(n4129)
         );
  OAI22_X1 U1017 ( .A1(n6749), .A2(n1702), .B1(n6747), .B2(n5781), .ZN(n4130)
         );
  BUF_X1 U1018 ( .A(n5096), .Z(n6274) );
  BUF_X1 U1019 ( .A(n5096), .Z(n6275) );
  BUF_X1 U1020 ( .A(n4397), .Z(n6488) );
  BUF_X1 U1021 ( .A(n4397), .Z(n6489) );
  NAND2_X1 U1022 ( .A1(n5730), .A2(n5736), .ZN(n6173) );
  NAND2_X1 U1023 ( .A1(n5730), .A2(n5736), .ZN(n5128) );
  NAND2_X1 U1024 ( .A1(n2893), .A2(n1786), .ZN(n2896) );
  NAND2_X1 U1025 ( .A1(n2893), .A2(n1750), .ZN(n2861) );
  NAND2_X1 U1026 ( .A1(n2616), .A2(n1786), .ZN(n2619) );
  NAND2_X1 U1027 ( .A1(n2616), .A2(n1750), .ZN(n2584) );
  NAND2_X1 U1028 ( .A1(n1894), .A2(n1786), .ZN(n1897) );
  NAND2_X1 U1029 ( .A1(n1894), .A2(n1750), .ZN(n1862) );
  NAND2_X1 U1030 ( .A1(n4319), .A2(n1786), .ZN(n4320) );
  NAND2_X1 U1031 ( .A1(n4319), .A2(n1750), .ZN(n4285) );
  NAND2_X1 U1032 ( .A1(n4182), .A2(n1786), .ZN(n4183) );
  NAND2_X1 U1033 ( .A1(n4182), .A2(n1750), .ZN(n4148) );
  NAND2_X1 U1034 ( .A1(n2755), .A2(n1786), .ZN(n2756) );
  NAND2_X1 U1035 ( .A1(n2755), .A2(n1750), .ZN(n2721) );
  NAND2_X1 U1036 ( .A1(n2031), .A2(n1786), .ZN(n2032) );
  NAND2_X1 U1037 ( .A1(n2031), .A2(n1750), .ZN(n1997) );
  BUF_X1 U1038 ( .A(n5096), .Z(n6276) );
  BUF_X1 U1039 ( .A(n4397), .Z(n6490) );
  NAND2_X1 U1040 ( .A1(n4319), .A2(n1856), .ZN(n4391) );
  NAND2_X1 U1041 ( .A1(n2893), .A2(n1856), .ZN(n2973) );
  NAND2_X1 U1042 ( .A1(n2616), .A2(n1856), .ZN(n2687) );
  NAND2_X1 U1043 ( .A1(n4182), .A2(n1856), .ZN(n4251) );
  NAND2_X1 U1044 ( .A1(n2755), .A2(n1856), .ZN(n2824) );
  NAND2_X1 U1045 ( .A1(n2031), .A2(n1856), .ZN(n2100) );
  NAND2_X1 U1046 ( .A1(n4319), .A2(n1821), .ZN(n4357) );
  NAND2_X1 U1047 ( .A1(n2893), .A2(n1821), .ZN(n2930) );
  NAND2_X1 U1048 ( .A1(n2616), .A2(n1821), .ZN(n2653) );
  NAND2_X1 U1049 ( .A1(n4182), .A2(n1821), .ZN(n4217) );
  NAND2_X1 U1050 ( .A1(n2755), .A2(n1821), .ZN(n2790) );
  NAND2_X1 U1051 ( .A1(n2031), .A2(n1821), .ZN(n2066) );
  AND3_X1 U1052 ( .A1(n1857), .A2(n1858), .A3(n2858), .ZN(n2755) );
  AND2_X1 U1053 ( .A1(n5725), .A2(n5738), .ZN(n5130) );
  NAND2_X1 U1054 ( .A1(n1894), .A2(n1856), .ZN(n6699) );
  NAND2_X1 U1055 ( .A1(n1894), .A2(n1856), .ZN(n1965) );
  NAND2_X1 U1056 ( .A1(n1894), .A2(n1821), .ZN(n6706) );
  NAND2_X1 U1057 ( .A1(n1894), .A2(n1821), .ZN(n1931) );
  AND2_X1 U1058 ( .A1(n5738), .A2(n5730), .ZN(n5125) );
  AND2_X1 U1059 ( .A1(n5727), .A2(n5730), .ZN(n5106) );
  AND2_X1 U1060 ( .A1(n5727), .A2(n5737), .ZN(n5135) );
  AND2_X1 U1061 ( .A1(n5733), .A2(n5727), .ZN(n5111) );
  AND2_X1 U1062 ( .A1(n5732), .A2(n5727), .ZN(n5112) );
  AND2_X1 U1063 ( .A1(n5733), .A2(n5738), .ZN(n5140) );
  AND2_X1 U1064 ( .A1(n5732), .A2(n5738), .ZN(n5141) );
  AND2_X1 U1065 ( .A1(n5726), .A2(n5738), .ZN(n5131) );
  AND2_X1 U1066 ( .A1(n5727), .A2(n5729), .ZN(n5107) );
  AND2_X1 U1067 ( .A1(n5738), .A2(n5729), .ZN(n5126) );
  AND2_X1 U1068 ( .A1(n5727), .A2(n5735), .ZN(n5136) );
  NOR3_X1 U1069 ( .A1(n5748), .A2(add_rd1[0]), .A3(n5744), .ZN(n5735) );
  NOR3_X1 U1070 ( .A1(n5744), .A2(add_rd1[4]), .A3(n5745), .ZN(n5730) );
  NOR2_X1 U1071 ( .A1(n5749), .A2(add_rd1[1]), .ZN(n5727) );
  NOR3_X1 U1072 ( .A1(n5748), .A2(add_rd1[3]), .A3(n5745), .ZN(n5733) );
  NOR3_X1 U1073 ( .A1(add_rd1[0]), .A2(add_rd1[3]), .A3(n5748), .ZN(n5732) );
  NAND2_X1 U1074 ( .A1(n5752), .A2(enable), .ZN(n6074) );
  NAND2_X1 U1075 ( .A1(n5752), .A2(enable), .ZN(n6075) );
  NAND2_X1 U1076 ( .A1(n5084), .A2(enable), .ZN(n6279) );
  NAND2_X1 U1077 ( .A1(n5084), .A2(enable), .ZN(n6280) );
  AND2_X1 U1078 ( .A1(add_wr[1]), .A2(add_wr[0]), .ZN(n1856) );
  AND2_X1 U1079 ( .A1(add_wr[1]), .A2(n4354), .ZN(n1821) );
  NAND2_X1 U1080 ( .A1(n5752), .A2(enable), .ZN(n5092) );
  NAND2_X1 U1081 ( .A1(n5084), .A2(enable), .ZN(n4393) );
  NOR3_X1 U1082 ( .A1(n2719), .A2(add_wr[4]), .A3(n2720), .ZN(n1859) );
  AOI221_X1 U1083 ( .B1(n6261), .B2(\registers[5][0] ), .C1(n6263), .C2(
        \registers[4][0] ), .A(n5723), .ZN(n5722) );
  OAI22_X1 U1084 ( .A1(n2561), .A2(n6266), .B1(n4288), .B2(n6272), .ZN(n5723)
         );
  AOI221_X1 U1085 ( .B1(n6262), .B2(\registers[5][1] ), .C1(n6264), .C2(
        \registers[4][1] ), .A(n5703), .ZN(n5702) );
  OAI22_X1 U1086 ( .A1(n2562), .A2(n6267), .B1(n4289), .B2(n6273), .ZN(n5703)
         );
  AOI221_X1 U1087 ( .B1(n6164), .B2(\registers[15][2] ), .C1(n6170), .C2(
        \registers[14][2] ), .A(n5692), .ZN(n5691) );
  OAI22_X1 U1088 ( .A1(n2771), .A2(n6174), .B1(n5764), .B2(n5129), .ZN(n5692)
         );
  AOI221_X1 U1089 ( .B1(n6261), .B2(\registers[5][3] ), .C1(n6263), .C2(
        \registers[4][3] ), .A(n5665), .ZN(n5664) );
  OAI22_X1 U1090 ( .A1(n2563), .A2(n6267), .B1(n4290), .B2(n6272), .ZN(n5665)
         );
  AOI221_X1 U1091 ( .B1(n6166), .B2(\registers[15][5] ), .C1(n6171), .C2(
        \registers[14][5] ), .A(n5635), .ZN(n5634) );
  OAI22_X1 U1092 ( .A1(n2772), .A2(n6177), .B1(n5765), .B2(n5129), .ZN(n5635)
         );
  AOI221_X1 U1093 ( .B1(n6167), .B2(\registers[15][8] ), .C1(n6172), .C2(
        \registers[14][8] ), .A(n5578), .ZN(n5577) );
  OAI22_X1 U1094 ( .A1(n2773), .A2(n6178), .B1(n5766), .B2(n5129), .ZN(n5578)
         );
  AOI221_X1 U1095 ( .B1(n6262), .B2(\registers[5][10] ), .C1(n6264), .C2(
        \registers[4][10] ), .A(n5532), .ZN(n5531) );
  OAI22_X1 U1096 ( .A1(n2564), .A2(n6266), .B1(n4291), .B2(n6273), .ZN(n5532)
         );
  AOI221_X1 U1097 ( .B1(n6167), .B2(\registers[15][11] ), .C1(n6170), .C2(
        \registers[14][11] ), .A(n5521), .ZN(n5520) );
  OAI22_X1 U1098 ( .A1(n2774), .A2(n6175), .B1(n5767), .B2(n5129), .ZN(n5521)
         );
  AOI221_X1 U1099 ( .B1(n6166), .B2(\registers[15][14] ), .C1(n6171), .C2(
        \registers[14][14] ), .A(n5464), .ZN(n5463) );
  OAI22_X1 U1100 ( .A1(n2775), .A2(n6176), .B1(n5768), .B2(n5129), .ZN(n5464)
         );
  AOI221_X1 U1101 ( .B1(n6168), .B2(\registers[15][17] ), .C1(n6172), .C2(
        \registers[14][17] ), .A(n5407), .ZN(n5406) );
  OAI22_X1 U1102 ( .A1(n2776), .A2(n6179), .B1(n5769), .B2(n5129), .ZN(n5407)
         );
  AOI221_X1 U1103 ( .B1(n6261), .B2(\registers[5][18] ), .C1(n6263), .C2(
        \registers[4][18] ), .A(n5380), .ZN(n5379) );
  OAI22_X1 U1104 ( .A1(n2565), .A2(n6266), .B1(n4292), .B2(n6272), .ZN(n5380)
         );
  AOI221_X1 U1105 ( .B1(n6262), .B2(\registers[5][19] ), .C1(n6264), .C2(
        \registers[4][19] ), .A(n5361), .ZN(n5360) );
  OAI22_X1 U1106 ( .A1(n2566), .A2(n6267), .B1(n4293), .B2(n6273), .ZN(n5361)
         );
  AOI221_X1 U1107 ( .B1(n6169), .B2(\registers[15][20] ), .C1(n6170), .C2(
        \registers[14][20] ), .A(n5350), .ZN(n5349) );
  OAI22_X1 U1108 ( .A1(n2777), .A2(n6174), .B1(n5770), .B2(n5129), .ZN(n5350)
         );
  AOI221_X1 U1109 ( .B1(n6261), .B2(\registers[5][21] ), .C1(n6263), .C2(
        \registers[4][21] ), .A(n5323), .ZN(n5322) );
  OAI22_X1 U1110 ( .A1(n2567), .A2(n6267), .B1(n4294), .B2(n6272), .ZN(n5323)
         );
  AOI221_X1 U1111 ( .B1(n6163), .B2(\registers[15][23] ), .C1(n6171), .C2(
        \registers[14][23] ), .A(n5293), .ZN(n5292) );
  OAI22_X1 U1112 ( .A1(n2778), .A2(n6177), .B1(n5771), .B2(n5129), .ZN(n5293)
         );
  AOI221_X1 U1113 ( .B1(n6164), .B2(\registers[15][26] ), .C1(n6172), .C2(
        \registers[14][26] ), .A(n5236), .ZN(n5235) );
  OAI22_X1 U1114 ( .A1(n2779), .A2(n6178), .B1(n5772), .B2(n5129), .ZN(n5236)
         );
  AOI221_X1 U1115 ( .B1(n6262), .B2(\registers[5][28] ), .C1(n6264), .C2(
        \registers[4][28] ), .A(n5190), .ZN(n5189) );
  OAI22_X1 U1116 ( .A1(n2568), .A2(n6266), .B1(n4295), .B2(n6273), .ZN(n5190)
         );
  AOI221_X1 U1117 ( .B1(n6165), .B2(\registers[15][29] ), .C1(n6170), .C2(
        \registers[14][29] ), .A(n5179), .ZN(n5178) );
  OAI22_X1 U1118 ( .A1(n2780), .A2(n6175), .B1(n5773), .B2(n5129), .ZN(n5179)
         );
  AOI221_X1 U1119 ( .B1(n6464), .B2(\registers[5][0] ), .C1(n6470), .C2(
        \registers[4][0] ), .A(n5055), .ZN(n5054) );
  OAI22_X1 U1120 ( .A1(n2561), .A2(n6474), .B1(n4288), .B2(n6482), .ZN(n5055)
         );
  AOI221_X1 U1121 ( .B1(n6465), .B2(\registers[5][1] ), .C1(n6471), .C2(
        \registers[4][1] ), .A(n5034), .ZN(n5033) );
  OAI22_X1 U1122 ( .A1(n2562), .A2(n6478), .B1(n4289), .B2(n6486), .ZN(n5034)
         );
  AOI221_X1 U1123 ( .B1(n6464), .B2(\registers[5][2] ), .C1(n4403), .C2(
        \registers[4][2] ), .A(n5014), .ZN(n5013) );
  OAI22_X1 U1124 ( .A1(n2781), .A2(n6478), .B1(n5774), .B2(n6481), .ZN(n5014)
         );
  AOI221_X1 U1125 ( .B1(n6465), .B2(\registers[5][3] ), .C1(n6470), .C2(
        \registers[4][3] ), .A(n4994), .ZN(n4993) );
  OAI22_X1 U1126 ( .A1(n2563), .A2(n6477), .B1(n4290), .B2(n6487), .ZN(n4994)
         );
  AOI221_X1 U1127 ( .B1(n6466), .B2(\registers[5][4] ), .C1(n6471), .C2(
        \registers[4][4] ), .A(n4974), .ZN(n4973) );
  OAI22_X1 U1128 ( .A1(n2754), .A2(n6473), .B1(n4347), .B2(n6481), .ZN(n4974)
         );
  AOI221_X1 U1129 ( .B1(n6467), .B2(\registers[5][5] ), .C1(n4403), .C2(
        \registers[4][5] ), .A(n4954), .ZN(n4953) );
  OAI22_X1 U1130 ( .A1(n2782), .A2(n6474), .B1(n5775), .B2(n6482), .ZN(n4954)
         );
  AOI221_X1 U1131 ( .B1(n6466), .B2(\registers[5][6] ), .C1(n6470), .C2(
        \registers[4][6] ), .A(n4934), .ZN(n4933) );
  OAI22_X1 U1132 ( .A1(n2758), .A2(n6475), .B1(n4348), .B2(n6483), .ZN(n4934)
         );
  AOI221_X1 U1133 ( .B1(n6467), .B2(\registers[5][7] ), .C1(n6471), .C2(
        \registers[4][7] ), .A(n4914), .ZN(n4913) );
  OAI22_X1 U1134 ( .A1(n2759), .A2(n6476), .B1(n4349), .B2(n6483), .ZN(n4914)
         );
  AOI221_X1 U1135 ( .B1(n6468), .B2(\registers[5][8] ), .C1(n4403), .C2(
        \registers[4][8] ), .A(n4894), .ZN(n4893) );
  OAI22_X1 U1136 ( .A1(n2783), .A2(n6475), .B1(n5776), .B2(n6484), .ZN(n4894)
         );
  AOI221_X1 U1137 ( .B1(n6469), .B2(\registers[5][9] ), .C1(n6470), .C2(
        \registers[4][9] ), .A(n4874), .ZN(n4873) );
  OAI22_X1 U1138 ( .A1(n2760), .A2(n6476), .B1(n4350), .B2(n6485), .ZN(n4874)
         );
  AOI221_X1 U1139 ( .B1(n6464), .B2(\registers[5][10] ), .C1(n6471), .C2(
        \registers[4][10] ), .A(n4854), .ZN(n4853) );
  OAI22_X1 U1140 ( .A1(n2564), .A2(n6477), .B1(n4291), .B2(n6486), .ZN(n4854)
         );
  AOI221_X1 U1141 ( .B1(n6465), .B2(\registers[5][11] ), .C1(n4403), .C2(
        \registers[4][11] ), .A(n4834), .ZN(n4833) );
  OAI22_X1 U1142 ( .A1(n2784), .A2(n6479), .B1(n5777), .B2(n6487), .ZN(n4834)
         );
  AOI221_X1 U1143 ( .B1(n6468), .B2(\registers[5][12] ), .C1(n6470), .C2(
        \registers[4][12] ), .A(n4814), .ZN(n4813) );
  OAI22_X1 U1144 ( .A1(n2761), .A2(n6473), .B1(n4351), .B2(n6481), .ZN(n4814)
         );
  AOI221_X1 U1145 ( .B1(n6469), .B2(\registers[5][13] ), .C1(n6471), .C2(
        \registers[4][13] ), .A(n4794), .ZN(n4793) );
  OAI22_X1 U1146 ( .A1(n2762), .A2(n6474), .B1(n4352), .B2(n6482), .ZN(n4794)
         );
  AOI221_X1 U1147 ( .B1(n6466), .B2(\registers[5][14] ), .C1(n4403), .C2(
        \registers[4][14] ), .A(n4774), .ZN(n4773) );
  OAI22_X1 U1148 ( .A1(n2785), .A2(n6475), .B1(n5778), .B2(n6482), .ZN(n4774)
         );
  AOI221_X1 U1149 ( .B1(n6467), .B2(\registers[5][15] ), .C1(n6470), .C2(
        \registers[4][15] ), .A(n4754), .ZN(n4753) );
  OAI22_X1 U1150 ( .A1(n2763), .A2(n6476), .B1(n4353), .B2(n6483), .ZN(n4754)
         );
  AOI221_X1 U1151 ( .B1(n6468), .B2(\registers[5][16] ), .C1(n6471), .C2(
        \registers[4][16] ), .A(n4734), .ZN(n4733) );
  OAI22_X1 U1152 ( .A1(n2764), .A2(n6474), .B1(n4356), .B2(n6484), .ZN(n4734)
         );
  AOI221_X1 U1153 ( .B1(n6469), .B2(\registers[5][17] ), .C1(n4403), .C2(
        \registers[4][17] ), .A(n4714), .ZN(n4713) );
  OAI22_X1 U1154 ( .A1(n2786), .A2(n6476), .B1(n5779), .B2(n6485), .ZN(n4714)
         );
  AOI221_X1 U1155 ( .B1(n6464), .B2(\registers[5][18] ), .C1(n6470), .C2(
        \registers[4][18] ), .A(n4694), .ZN(n4693) );
  OAI22_X1 U1156 ( .A1(n2565), .A2(n6477), .B1(n4292), .B2(n6486), .ZN(n4694)
         );
  AOI221_X1 U1157 ( .B1(n6465), .B2(\registers[5][19] ), .C1(n6471), .C2(
        \registers[4][19] ), .A(n4674), .ZN(n4673) );
  OAI22_X1 U1158 ( .A1(n2566), .A2(n6478), .B1(n4293), .B2(n6487), .ZN(n4674)
         );
  AOI221_X1 U1159 ( .B1(n6464), .B2(\registers[5][20] ), .C1(n4403), .C2(
        \registers[4][20] ), .A(n4654), .ZN(n4653) );
  OAI22_X1 U1160 ( .A1(n2787), .A2(n6478), .B1(n5780), .B2(n6481), .ZN(n4654)
         );
  AOI221_X1 U1161 ( .B1(n6465), .B2(\registers[5][21] ), .C1(n6470), .C2(
        \registers[4][21] ), .A(n4634), .ZN(n4633) );
  OAI22_X1 U1162 ( .A1(n2567), .A2(n6479), .B1(n4294), .B2(n6485), .ZN(n4634)
         );
  AOI221_X1 U1163 ( .B1(n6466), .B2(\registers[5][22] ), .C1(n6471), .C2(
        \registers[4][22] ), .A(n4614), .ZN(n4613) );
  OAI22_X1 U1164 ( .A1(n2765), .A2(n6473), .B1(n4390), .B2(n6487), .ZN(n4614)
         );
  AOI221_X1 U1165 ( .B1(n6467), .B2(\registers[5][23] ), .C1(n4403), .C2(
        \registers[4][23] ), .A(n4594), .ZN(n4593) );
  OAI22_X1 U1166 ( .A1(n2788), .A2(n6478), .B1(n5781), .B2(n6486), .ZN(n4594)
         );
  AOI221_X1 U1167 ( .B1(n6466), .B2(\registers[5][24] ), .C1(n6470), .C2(
        \registers[4][24] ), .A(n4574), .ZN(n4573) );
  OAI22_X1 U1168 ( .A1(n2766), .A2(n6477), .B1(n5759), .B2(n6485), .ZN(n4574)
         );
  AOI221_X1 U1169 ( .B1(n6467), .B2(\registers[5][25] ), .C1(n6471), .C2(
        \registers[4][25] ), .A(n4554), .ZN(n4553) );
  OAI22_X1 U1170 ( .A1(n2767), .A2(n6477), .B1(n5760), .B2(n6487), .ZN(n4554)
         );
  AOI221_X1 U1171 ( .B1(n6468), .B2(\registers[5][26] ), .C1(n4403), .C2(
        \registers[4][26] ), .A(n4534), .ZN(n4533) );
  OAI22_X1 U1172 ( .A1(n2789), .A2(n6473), .B1(n5782), .B2(n6484), .ZN(n4534)
         );
  AOI221_X1 U1173 ( .B1(n6469), .B2(\registers[5][27] ), .C1(n6470), .C2(
        \registers[4][27] ), .A(n4514), .ZN(n4513) );
  OAI22_X1 U1174 ( .A1(n2768), .A2(n6479), .B1(n5761), .B2(n6484), .ZN(n4514)
         );
  AOI221_X1 U1175 ( .B1(n6464), .B2(\registers[5][28] ), .C1(n6471), .C2(
        \registers[4][28] ), .A(n4494), .ZN(n4493) );
  OAI22_X1 U1176 ( .A1(n2568), .A2(n6475), .B1(n4295), .B2(n6483), .ZN(n4494)
         );
  AOI221_X1 U1177 ( .B1(n6465), .B2(\registers[5][29] ), .C1(n4403), .C2(
        \registers[4][29] ), .A(n4474), .ZN(n4473) );
  OAI22_X1 U1178 ( .A1(n2791), .A2(n6479), .B1(n5783), .B2(n6481), .ZN(n4474)
         );
  AOI221_X1 U1179 ( .B1(n6468), .B2(\registers[5][30] ), .C1(n6470), .C2(
        \registers[4][30] ), .A(n4454), .ZN(n4453) );
  OAI22_X1 U1180 ( .A1(n2769), .A2(n6479), .B1(n5762), .B2(n6486), .ZN(n4454)
         );
  AOI221_X1 U1181 ( .B1(n6469), .B2(\registers[5][31] ), .C1(n6471), .C2(
        \registers[4][31] ), .A(n4404), .ZN(n4401) );
  OAI22_X1 U1182 ( .A1(n2770), .A2(n6473), .B1(n5763), .B2(n6483), .ZN(n4404)
         );
  AOI221_X1 U1183 ( .B1(n6136), .B2(\registers[6][0] ), .C1(n6144), .C2(
        \registers[7][0] ), .A(n5746), .ZN(n5741) );
  OAI22_X1 U1184 ( .A1(n2569), .A2(n6152), .B1(n4296), .B2(n6159), .ZN(n5746)
         );
  AOI221_X1 U1185 ( .B1(n6142), .B2(\registers[6][1] ), .C1(n6145), .C2(
        \registers[7][1] ), .A(n5712), .ZN(n5709) );
  OAI22_X1 U1186 ( .A1(n2570), .A2(n6151), .B1(n4297), .B2(n6158), .ZN(n5712)
         );
  AOI221_X1 U1187 ( .B1(n6136), .B2(\registers[6][2] ), .C1(n6143), .C2(
        \registers[7][2] ), .A(n5693), .ZN(n5690) );
  OAI22_X1 U1188 ( .A1(n2571), .A2(n6151), .B1(n4298), .B2(n6159), .ZN(n5693)
         );
  AOI221_X1 U1189 ( .B1(n6138), .B2(\registers[6][3] ), .C1(n6143), .C2(
        \registers[7][3] ), .A(n5674), .ZN(n5671) );
  OAI22_X1 U1190 ( .A1(n2572), .A2(n6150), .B1(n4299), .B2(n6155), .ZN(n5674)
         );
  AOI221_X1 U1191 ( .B1(n6139), .B2(\registers[6][4] ), .C1(n6144), .C2(
        \registers[7][4] ), .A(n5655), .ZN(n5652) );
  OAI22_X1 U1192 ( .A1(n2573), .A2(n6147), .B1(n4300), .B2(n6155), .ZN(n5655)
         );
  AOI221_X1 U1193 ( .B1(n6136), .B2(\registers[6][5] ), .C1(n6144), .C2(
        \registers[7][5] ), .A(n5636), .ZN(n5633) );
  OAI22_X1 U1194 ( .A1(n2574), .A2(n6148), .B1(n4301), .B2(n6156), .ZN(n5636)
         );
  AOI221_X1 U1195 ( .B1(n6137), .B2(\registers[6][6] ), .C1(n6145), .C2(
        \registers[7][6] ), .A(n5617), .ZN(n5614) );
  OAI22_X1 U1196 ( .A1(n2575), .A2(n6149), .B1(n4302), .B2(n6157), .ZN(n5617)
         );
  AOI221_X1 U1197 ( .B1(n6138), .B2(\registers[6][7] ), .C1(n6143), .C2(
        \registers[7][7] ), .A(n5598), .ZN(n5595) );
  OAI22_X1 U1198 ( .A1(n2576), .A2(n6149), .B1(n4303), .B2(n6158), .ZN(n5598)
         );
  AOI221_X1 U1199 ( .B1(n6137), .B2(\registers[6][8] ), .C1(n6145), .C2(
        \registers[7][8] ), .A(n5579), .ZN(n5576) );
  OAI22_X1 U1200 ( .A1(n2577), .A2(n6150), .B1(n4304), .B2(n6156), .ZN(n5579)
         );
  AOI221_X1 U1201 ( .B1(n6140), .B2(\registers[6][9] ), .C1(n6144), .C2(
        \registers[7][9] ), .A(n5560), .ZN(n5557) );
  OAI22_X1 U1202 ( .A1(n2578), .A2(n6151), .B1(n4305), .B2(n6158), .ZN(n5560)
         );
  AOI221_X1 U1203 ( .B1(n6139), .B2(\registers[6][10] ), .C1(n6145), .C2(
        \registers[7][10] ), .A(n5541), .ZN(n5538) );
  OAI22_X1 U1204 ( .A1(n2579), .A2(n6152), .B1(n4306), .B2(n6159), .ZN(n5541)
         );
  AOI221_X1 U1205 ( .B1(n6140), .B2(\registers[6][11] ), .C1(n6143), .C2(
        \registers[7][11] ), .A(n5522), .ZN(n5519) );
  OAI22_X1 U1206 ( .A1(n2580), .A2(n6153), .B1(n4307), .B2(n6161), .ZN(n5522)
         );
  AOI221_X1 U1207 ( .B1(n6141), .B2(\registers[6][12] ), .C1(n6143), .C2(
        \registers[7][12] ), .A(n5503), .ZN(n5500) );
  OAI22_X1 U1208 ( .A1(n2581), .A2(n6147), .B1(n4308), .B2(n6155), .ZN(n5503)
         );
  AOI221_X1 U1209 ( .B1(n6141), .B2(\registers[6][13] ), .C1(n6144), .C2(
        \registers[7][13] ), .A(n5484), .ZN(n5481) );
  OAI22_X1 U1210 ( .A1(n2583), .A2(n6148), .B1(n4309), .B2(n6156), .ZN(n5484)
         );
  AOI221_X1 U1211 ( .B1(n6139), .B2(\registers[6][14] ), .C1(n6144), .C2(
        \registers[7][14] ), .A(n5465), .ZN(n5462) );
  OAI22_X1 U1212 ( .A1(n2618), .A2(n6149), .B1(n4310), .B2(n6157), .ZN(n5465)
         );
  AOI221_X1 U1213 ( .B1(n6140), .B2(\registers[6][15] ), .C1(n6145), .C2(
        \registers[7][15] ), .A(n5446), .ZN(n5443) );
  OAI22_X1 U1214 ( .A1(n2652), .A2(n6149), .B1(n4311), .B2(n6158), .ZN(n5446)
         );
  AOI221_X1 U1215 ( .B1(n6141), .B2(\registers[6][16] ), .C1(n6143), .C2(
        \registers[7][16] ), .A(n5427), .ZN(n5424) );
  OAI22_X1 U1216 ( .A1(n2686), .A2(n6150), .B1(n4312), .B2(n6157), .ZN(n5427)
         );
  AOI221_X1 U1217 ( .B1(n6141), .B2(\registers[6][17] ), .C1(n6145), .C2(
        \registers[7][17] ), .A(n5408), .ZN(n5405) );
  OAI22_X1 U1218 ( .A1(n2723), .A2(n6151), .B1(n4313), .B2(n6157), .ZN(n5408)
         );
  AOI221_X1 U1219 ( .B1(n6142), .B2(\registers[6][18] ), .C1(n6144), .C2(
        \registers[7][18] ), .A(n5389), .ZN(n5386) );
  OAI22_X1 U1220 ( .A1(n2724), .A2(n6152), .B1(n4314), .B2(n6159), .ZN(n5389)
         );
  AOI221_X1 U1221 ( .B1(n6142), .B2(\registers[6][19] ), .C1(n6145), .C2(
        \registers[7][19] ), .A(n5370), .ZN(n5367) );
  OAI22_X1 U1222 ( .A1(n2725), .A2(n6153), .B1(n4315), .B2(n6160), .ZN(n5370)
         );
  AOI221_X1 U1223 ( .B1(n6142), .B2(\registers[6][20] ), .C1(n6143), .C2(
        \registers[7][20] ), .A(n5351), .ZN(n5348) );
  OAI22_X1 U1224 ( .A1(n2726), .A2(n6153), .B1(n4316), .B2(n6160), .ZN(n5351)
         );
  AOI221_X1 U1225 ( .B1(n6142), .B2(\registers[6][21] ), .C1(n6143), .C2(
        \registers[7][21] ), .A(n5332), .ZN(n5329) );
  OAI22_X1 U1226 ( .A1(n2727), .A2(n6148), .B1(n4317), .B2(n6160), .ZN(n5332)
         );
  AOI221_X1 U1227 ( .B1(n6137), .B2(\registers[6][28] ), .C1(n6145), .C2(
        \registers[7][28] ), .A(n5199), .ZN(n5196) );
  OAI22_X1 U1228 ( .A1(n2728), .A2(n6153), .B1(n4318), .B2(n6161), .ZN(n5199)
         );
  AOI221_X1 U1229 ( .B1(n6138), .B2(\registers[6][29] ), .C1(n6143), .C2(
        \registers[7][29] ), .A(n5180), .ZN(n5177) );
  OAI22_X1 U1230 ( .A1(n2729), .A2(n6150), .B1(n4322), .B2(n6156), .ZN(n5180)
         );
  AOI221_X1 U1231 ( .B1(n6138), .B2(\registers[6][30] ), .C1(n6143), .C2(
        \registers[7][30] ), .A(n5161), .ZN(n5158) );
  OAI22_X1 U1232 ( .A1(n2730), .A2(n6148), .B1(n4323), .B2(n6160), .ZN(n5161)
         );
  AOI221_X1 U1233 ( .B1(n6139), .B2(\registers[6][31] ), .C1(n6144), .C2(
        \registers[7][31] ), .A(n5132), .ZN(n5123) );
  OAI22_X1 U1234 ( .A1(n2731), .A2(n6148), .B1(n4324), .B2(n6161), .ZN(n5132)
         );
  AOI221_X1 U1235 ( .B1(n6432), .B2(\registers[13][0] ), .C1(n6440), .C2(
        \registers[12][0] ), .A(n5060), .ZN(n5053) );
  OAI22_X1 U1236 ( .A1(n2792), .A2(n6451), .B1(n5784), .B2(n6460), .ZN(n5060)
         );
  AOI221_X1 U1237 ( .B1(n6341), .B2(\registers[6][0] ), .C1(n6348), .C2(
        \registers[7][0] ), .A(n5078), .ZN(n5073) );
  OAI22_X1 U1238 ( .A1(n2569), .A2(n6359), .B1(n4296), .B2(n6368), .ZN(n5078)
         );
  AOI221_X1 U1239 ( .B1(n6433), .B2(\registers[13][1] ), .C1(n6440), .C2(
        \registers[12][1] ), .A(n5035), .ZN(n5032) );
  OAI22_X1 U1240 ( .A1(n2794), .A2(n6453), .B1(n5786), .B2(n6462), .ZN(n5035)
         );
  AOI221_X1 U1241 ( .B1(n6345), .B2(\registers[6][1] ), .C1(n6348), .C2(
        \registers[7][1] ), .A(n5043), .ZN(n5040) );
  OAI22_X1 U1242 ( .A1(n2570), .A2(n6362), .B1(n4297), .B2(n6364), .ZN(n5043)
         );
  AOI221_X1 U1243 ( .B1(n6432), .B2(\registers[13][2] ), .C1(n6444), .C2(
        \registers[12][2] ), .A(n5015), .ZN(n5012) );
  OAI22_X1 U1244 ( .A1(n2796), .A2(n6454), .B1(n5788), .B2(n6461), .ZN(n5015)
         );
  AOI221_X1 U1245 ( .B1(n6341), .B2(\registers[6][2] ), .C1(n6349), .C2(
        \registers[7][2] ), .A(n5023), .ZN(n5020) );
  OAI22_X1 U1246 ( .A1(n2571), .A2(n6360), .B1(n4298), .B2(n6369), .ZN(n5023)
         );
  AOI221_X1 U1247 ( .B1(n6432), .B2(\registers[13][3] ), .C1(n6441), .C2(
        \registers[12][3] ), .A(n4995), .ZN(n4992) );
  OAI22_X1 U1248 ( .A1(n2798), .A2(n6452), .B1(n5790), .B2(n6460), .ZN(n4995)
         );
  AOI221_X1 U1249 ( .B1(n6342), .B2(\registers[6][3] ), .C1(n6351), .C2(
        \registers[7][3] ), .A(n5003), .ZN(n5000) );
  OAI22_X1 U1250 ( .A1(n2572), .A2(n6357), .B1(n4299), .B2(n6369), .ZN(n5003)
         );
  AOI221_X1 U1251 ( .B1(n6435), .B2(\registers[13][4] ), .C1(n6442), .C2(
        \registers[12][4] ), .A(n4975), .ZN(n4972) );
  OAI22_X1 U1252 ( .A1(n2800), .A2(n6448), .B1(n5792), .B2(n6456), .ZN(n4975)
         );
  AOI221_X1 U1253 ( .B1(n6343), .B2(\registers[6][4] ), .C1(n6348), .C2(
        \registers[7][4] ), .A(n4983), .ZN(n4980) );
  OAI22_X1 U1254 ( .A1(n2573), .A2(n6356), .B1(n4300), .B2(n6364), .ZN(n4983)
         );
  AOI221_X1 U1255 ( .B1(n6432), .B2(\registers[13][5] ), .C1(n6441), .C2(
        \registers[12][5] ), .A(n4955), .ZN(n4952) );
  OAI22_X1 U1256 ( .A1(n2802), .A2(n6449), .B1(n5794), .B2(n6457), .ZN(n4955)
         );
  AOI221_X1 U1257 ( .B1(n6342), .B2(\registers[6][5] ), .C1(n6348), .C2(
        \registers[7][5] ), .A(n4963), .ZN(n4960) );
  OAI22_X1 U1258 ( .A1(n2574), .A2(n6357), .B1(n4301), .B2(n6365), .ZN(n4963)
         );
  AOI221_X1 U1259 ( .B1(n6434), .B2(\registers[13][6] ), .C1(n6443), .C2(
        \registers[12][6] ), .A(n4935), .ZN(n4932) );
  OAI22_X1 U1260 ( .A1(n2804), .A2(n6450), .B1(n5796), .B2(n6458), .ZN(n4935)
         );
  AOI221_X1 U1261 ( .B1(n6344), .B2(\registers[6][6] ), .C1(n6350), .C2(
        \registers[7][6] ), .A(n4943), .ZN(n4940) );
  OAI22_X1 U1262 ( .A1(n2575), .A2(n6358), .B1(n4302), .B2(n6366), .ZN(n4943)
         );
  AOI221_X1 U1263 ( .B1(n6436), .B2(\registers[13][7] ), .C1(n6446), .C2(
        \registers[12][7] ), .A(n4915), .ZN(n4912) );
  OAI22_X1 U1264 ( .A1(n2806), .A2(n6451), .B1(n5798), .B2(n6457), .ZN(n4915)
         );
  AOI221_X1 U1265 ( .B1(n6346), .B2(\registers[6][7] ), .C1(n6352), .C2(
        \registers[7][7] ), .A(n4923), .ZN(n4920) );
  OAI22_X1 U1266 ( .A1(n2576), .A2(n6358), .B1(n4303), .B2(n6367), .ZN(n4923)
         );
  AOI221_X1 U1267 ( .B1(n6434), .B2(\registers[13][8] ), .C1(n6443), .C2(
        \registers[12][8] ), .A(n4895), .ZN(n4892) );
  OAI22_X1 U1268 ( .A1(n2808), .A2(n6451), .B1(n5800), .B2(n6457), .ZN(n4895)
         );
  AOI221_X1 U1269 ( .B1(n6343), .B2(\registers[6][8] ), .C1(n6350), .C2(
        \registers[7][8] ), .A(n4903), .ZN(n4900) );
  OAI22_X1 U1270 ( .A1(n2577), .A2(n6359), .B1(n4304), .B2(n6367), .ZN(n4903)
         );
  AOI221_X1 U1271 ( .B1(n6436), .B2(\registers[13][9] ), .C1(n6444), .C2(
        \registers[12][9] ), .A(n4875), .ZN(n4872) );
  OAI22_X1 U1272 ( .A1(n2810), .A2(n6449), .B1(n5802), .B2(n6459), .ZN(n4875)
         );
  AOI221_X1 U1273 ( .B1(n6344), .B2(\registers[6][9] ), .C1(n6352), .C2(
        \registers[7][9] ), .A(n4883), .ZN(n4880) );
  OAI22_X1 U1274 ( .A1(n2578), .A2(n6360), .B1(n4305), .B2(n6366), .ZN(n4883)
         );
  AOI221_X1 U1275 ( .B1(n6435), .B2(\registers[13][10] ), .C1(n6444), .C2(
        \registers[12][10] ), .A(n4855), .ZN(n4852) );
  OAI22_X1 U1276 ( .A1(n2812), .A2(n6452), .B1(n5804), .B2(n6456), .ZN(n4855)
         );
  AOI221_X1 U1277 ( .B1(n6343), .B2(\registers[6][10] ), .C1(n6351), .C2(
        \registers[7][10] ), .A(n4863), .ZN(n4860) );
  OAI22_X1 U1278 ( .A1(n2579), .A2(n6361), .B1(n4306), .B2(n6364), .ZN(n4863)
         );
  AOI221_X1 U1279 ( .B1(n6436), .B2(\registers[13][11] ), .C1(n6442), .C2(
        \registers[12][11] ), .A(n4835), .ZN(n4832) );
  OAI22_X1 U1280 ( .A1(n2814), .A2(n6453), .B1(n5806), .B2(n6460), .ZN(n4835)
         );
  AOI221_X1 U1281 ( .B1(n6344), .B2(\registers[6][11] ), .C1(n6352), .C2(
        \registers[7][11] ), .A(n4843), .ZN(n4840) );
  OAI22_X1 U1282 ( .A1(n2580), .A2(n6361), .B1(n4307), .B2(n6368), .ZN(n4843)
         );
  AOI221_X1 U1283 ( .B1(n6437), .B2(\registers[13][12] ), .C1(n6445), .C2(
        \registers[12][12] ), .A(n4815), .ZN(n4812) );
  OAI22_X1 U1284 ( .A1(n2816), .A2(n6448), .B1(n5808), .B2(n6456), .ZN(n4815)
         );
  AOI221_X1 U1285 ( .B1(n6345), .B2(\registers[6][12] ), .C1(n6353), .C2(
        \registers[7][12] ), .A(n4823), .ZN(n4820) );
  OAI22_X1 U1286 ( .A1(n2581), .A2(n6356), .B1(n4308), .B2(n6364), .ZN(n4823)
         );
  AOI221_X1 U1287 ( .B1(n6437), .B2(\registers[13][13] ), .C1(n6445), .C2(
        \registers[12][13] ), .A(n4795), .ZN(n4792) );
  OAI22_X1 U1288 ( .A1(n2818), .A2(n6449), .B1(n5810), .B2(n6457), .ZN(n4795)
         );
  AOI221_X1 U1289 ( .B1(n6345), .B2(\registers[6][13] ), .C1(n6353), .C2(
        \registers[7][13] ), .A(n4803), .ZN(n4800) );
  OAI22_X1 U1290 ( .A1(n2583), .A2(n6357), .B1(n4309), .B2(n6365), .ZN(n4803)
         );
  AOI221_X1 U1291 ( .B1(n6435), .B2(\registers[13][14] ), .C1(n6444), .C2(
        \registers[12][14] ), .A(n4775), .ZN(n4772) );
  OAI22_X1 U1292 ( .A1(n2820), .A2(n6450), .B1(n5812), .B2(n6458), .ZN(n4775)
         );
  AOI221_X1 U1293 ( .B1(n6343), .B2(\registers[6][14] ), .C1(n6351), .C2(
        \registers[7][14] ), .A(n4783), .ZN(n4780) );
  OAI22_X1 U1294 ( .A1(n2618), .A2(n6358), .B1(n4310), .B2(n6366), .ZN(n4783)
         );
  AOI221_X1 U1295 ( .B1(n6436), .B2(\registers[13][15] ), .C1(n6445), .C2(
        \registers[12][15] ), .A(n4755), .ZN(n4752) );
  OAI22_X1 U1296 ( .A1(n2822), .A2(n6451), .B1(n5814), .B2(n6459), .ZN(n4755)
         );
  AOI221_X1 U1297 ( .B1(n6344), .B2(\registers[6][15] ), .C1(n6352), .C2(
        \registers[7][15] ), .A(n4763), .ZN(n4760) );
  OAI22_X1 U1298 ( .A1(n2652), .A2(n6358), .B1(n4311), .B2(n6367), .ZN(n4763)
         );
  AOI221_X1 U1299 ( .B1(n6437), .B2(\registers[13][16] ), .C1(n6444), .C2(
        \registers[12][16] ), .A(n4735), .ZN(n4732) );
  OAI22_X1 U1300 ( .A1(n2826), .A2(n6449), .B1(n5816), .B2(n6459), .ZN(n4735)
         );
  AOI221_X1 U1301 ( .B1(n6345), .B2(\registers[6][16] ), .C1(n6353), .C2(
        \registers[7][16] ), .A(n4743), .ZN(n4740) );
  OAI22_X1 U1302 ( .A1(n2686), .A2(n6359), .B1(n4312), .B2(n6365), .ZN(n4743)
         );
  AOI221_X1 U1303 ( .B1(n6437), .B2(\registers[13][17] ), .C1(n6445), .C2(
        \registers[12][17] ), .A(n4715), .ZN(n4712) );
  OAI22_X1 U1304 ( .A1(n2828), .A2(n6450), .B1(n5818), .B2(n6459), .ZN(n4715)
         );
  AOI221_X1 U1305 ( .B1(n6345), .B2(\registers[6][17] ), .C1(n6353), .C2(
        \registers[7][17] ), .A(n4723), .ZN(n4720) );
  OAI22_X1 U1306 ( .A1(n2723), .A2(n6360), .B1(n4313), .B2(n6366), .ZN(n4723)
         );
  AOI221_X1 U1307 ( .B1(n6438), .B2(\registers[13][18] ), .C1(n6445), .C2(
        \registers[12][18] ), .A(n4695), .ZN(n4692) );
  OAI22_X1 U1308 ( .A1(n2830), .A2(n6452), .B1(n5820), .B2(n6461), .ZN(n4695)
         );
  AOI221_X1 U1309 ( .B1(n6346), .B2(\registers[6][18] ), .C1(n6354), .C2(
        \registers[7][18] ), .A(n4703), .ZN(n4700) );
  OAI22_X1 U1310 ( .A1(n2724), .A2(n6361), .B1(n4314), .B2(n6370), .ZN(n4703)
         );
  AOI221_X1 U1311 ( .B1(n6438), .B2(\registers[13][19] ), .C1(n6446), .C2(
        \registers[12][19] ), .A(n4675), .ZN(n4672) );
  OAI22_X1 U1312 ( .A1(n2832), .A2(n6453), .B1(n5822), .B2(n6462), .ZN(n4675)
         );
  AOI221_X1 U1313 ( .B1(n6346), .B2(\registers[6][19] ), .C1(n6354), .C2(
        \registers[7][19] ), .A(n4683), .ZN(n4680) );
  OAI22_X1 U1314 ( .A1(n2725), .A2(n6361), .B1(n4315), .B2(n6368), .ZN(n4683)
         );
  AOI221_X1 U1315 ( .B1(n6438), .B2(\registers[13][20] ), .C1(n6446), .C2(
        \registers[12][20] ), .A(n4655), .ZN(n4652) );
  OAI22_X1 U1316 ( .A1(n2834), .A2(n6454), .B1(n5824), .B2(n6460), .ZN(n4655)
         );
  AOI221_X1 U1317 ( .B1(n6346), .B2(\registers[6][20] ), .C1(n6354), .C2(
        \registers[7][20] ), .A(n4663), .ZN(n4660) );
  OAI22_X1 U1318 ( .A1(n2726), .A2(n6362), .B1(n4316), .B2(n6369), .ZN(n4663)
         );
  AOI221_X1 U1319 ( .B1(n6438), .B2(\registers[13][21] ), .C1(n6446), .C2(
        \registers[12][21] ), .A(n4635), .ZN(n4632) );
  OAI22_X1 U1320 ( .A1(n2836), .A2(n6452), .B1(n5826), .B2(n6460), .ZN(n4635)
         );
  AOI221_X1 U1321 ( .B1(n6346), .B2(\registers[6][21] ), .C1(n6354), .C2(
        \registers[7][21] ), .A(n4643), .ZN(n4640) );
  OAI22_X1 U1322 ( .A1(n2727), .A2(n6357), .B1(n4317), .B2(n6369), .ZN(n4643)
         );
  AOI221_X1 U1323 ( .B1(n6432), .B2(\registers[13][22] ), .C1(n6440), .C2(
        \registers[12][22] ), .A(n4615), .ZN(n4612) );
  OAI22_X1 U1324 ( .A1(n2838), .A2(n6454), .B1(n5828), .B2(n6461), .ZN(n4615)
         );
  AOI221_X1 U1325 ( .B1(n6341), .B2(\registers[6][22] ), .C1(n6348), .C2(
        \registers[7][22] ), .A(n4623), .ZN(n4620) );
  OAI22_X1 U1326 ( .A1(n4202), .A2(n6361), .B1(n5901), .B2(n6370), .ZN(n4623)
         );
  AOI221_X1 U1327 ( .B1(n6433), .B2(\registers[13][23] ), .C1(n6440), .C2(
        \registers[12][23] ), .A(n4595), .ZN(n4592) );
  OAI22_X1 U1328 ( .A1(n2839), .A2(n6448), .B1(n5829), .B2(n6462), .ZN(n4595)
         );
  AOI221_X1 U1329 ( .B1(n6345), .B2(\registers[6][23] ), .C1(n6349), .C2(
        \registers[7][23] ), .A(n4603), .ZN(n4600) );
  OAI22_X1 U1330 ( .A1(n4204), .A2(n6362), .B1(n5903), .B2(n6368), .ZN(n4603)
         );
  AOI221_X1 U1331 ( .B1(n6433), .B2(\registers[13][24] ), .C1(n6440), .C2(
        \registers[12][24] ), .A(n4575), .ZN(n4572) );
  OAI22_X1 U1332 ( .A1(n2840), .A2(n6453), .B1(n5830), .B2(n6458), .ZN(n4575)
         );
  AOI221_X1 U1333 ( .B1(n6346), .B2(\registers[6][24] ), .C1(n6349), .C2(
        \registers[7][24] ), .A(n4583), .ZN(n4580) );
  OAI22_X1 U1334 ( .A1(n4206), .A2(n6356), .B1(n5905), .B2(n6367), .ZN(n4583)
         );
  AOI221_X1 U1335 ( .B1(n6437), .B2(\registers[13][25] ), .C1(n6441), .C2(
        \registers[12][25] ), .A(n4555), .ZN(n4552) );
  OAI22_X1 U1336 ( .A1(n2841), .A2(n6454), .B1(n5831), .B2(n6462), .ZN(n4555)
         );
  AOI221_X1 U1337 ( .B1(n6342), .B2(\registers[6][25] ), .C1(n6352), .C2(
        \registers[7][25] ), .A(n4563), .ZN(n4560) );
  OAI22_X1 U1338 ( .A1(n4208), .A2(n6362), .B1(n5907), .B2(n6369), .ZN(n4563)
         );
  AOI221_X1 U1339 ( .B1(n6434), .B2(\registers[13][26] ), .C1(n6442), .C2(
        \registers[12][26] ), .A(n4535), .ZN(n4532) );
  OAI22_X1 U1340 ( .A1(n2842), .A2(n6452), .B1(n5832), .B2(n6458), .ZN(n4535)
         );
  AOI221_X1 U1341 ( .B1(n6343), .B2(\registers[6][26] ), .C1(n6351), .C2(
        \registers[7][26] ), .A(n4543), .ZN(n4540) );
  OAI22_X1 U1342 ( .A1(n4210), .A2(n6362), .B1(n5909), .B2(n6365), .ZN(n4543)
         );
  AOI221_X1 U1343 ( .B1(n6435), .B2(\registers[13][27] ), .C1(n6442), .C2(
        \registers[12][27] ), .A(n4515), .ZN(n4512) );
  OAI22_X1 U1344 ( .A1(n2843), .A2(n6453), .B1(n5833), .B2(n6461), .ZN(n4515)
         );
  AOI221_X1 U1345 ( .B1(n6342), .B2(\registers[6][27] ), .C1(n6353), .C2(
        \registers[7][27] ), .A(n4523), .ZN(n4520) );
  OAI22_X1 U1346 ( .A1(n4212), .A2(n6356), .B1(n5911), .B2(n6370), .ZN(n4523)
         );
  AOI221_X1 U1347 ( .B1(n6434), .B2(\registers[13][28] ), .C1(n6443), .C2(
        \registers[12][28] ), .A(n4495), .ZN(n4492) );
  OAI22_X1 U1348 ( .A1(n2844), .A2(n6450), .B1(n5834), .B2(n6456), .ZN(n4495)
         );
  AOI221_X1 U1349 ( .B1(n6341), .B2(\registers[6][28] ), .C1(n6350), .C2(
        \registers[7][28] ), .A(n4503), .ZN(n4500) );
  OAI22_X1 U1350 ( .A1(n2728), .A2(n6360), .B1(n4318), .B2(n6364), .ZN(n4503)
         );
  AOI221_X1 U1351 ( .B1(n6434), .B2(\registers[13][29] ), .C1(n6446), .C2(
        \registers[12][29] ), .A(n4475), .ZN(n4472) );
  OAI22_X1 U1352 ( .A1(n2846), .A2(n6454), .B1(n5836), .B2(n6461), .ZN(n4475)
         );
  AOI221_X1 U1353 ( .B1(n6341), .B2(\registers[6][29] ), .C1(n6350), .C2(
        \registers[7][29] ), .A(n4483), .ZN(n4480) );
  OAI22_X1 U1354 ( .A1(n2729), .A2(n6356), .B1(n4322), .B2(n6370), .ZN(n4483)
         );
  AOI221_X1 U1355 ( .B1(n6433), .B2(\registers[13][30] ), .C1(n6441), .C2(
        \registers[12][30] ), .A(n4455), .ZN(n4452) );
  OAI22_X1 U1356 ( .A1(n2848), .A2(n6448), .B1(n5838), .B2(n6456), .ZN(n4455)
         );
  AOI221_X1 U1357 ( .B1(n6344), .B2(\registers[6][30] ), .C1(n6349), .C2(
        \registers[7][30] ), .A(n4463), .ZN(n4460) );
  OAI22_X1 U1358 ( .A1(n2730), .A2(n6357), .B1(n4323), .B2(n6370), .ZN(n4463)
         );
  AOI221_X1 U1359 ( .B1(n6435), .B2(\registers[13][31] ), .C1(n6443), .C2(
        \registers[12][31] ), .A(n4409), .ZN(n4400) );
  OAI22_X1 U1360 ( .A1(n2850), .A2(n6448), .B1(n5840), .B2(n6462), .ZN(n4409)
         );
  AOI221_X1 U1361 ( .B1(n6343), .B2(\registers[6][31] ), .C1(n6351), .C2(
        \registers[7][31] ), .A(n4433), .ZN(n4424) );
  OAI22_X1 U1362 ( .A1(n2731), .A2(n6359), .B1(n4324), .B2(n6368), .ZN(n4433)
         );
  AOI221_X1 U1363 ( .B1(n6168), .B2(\registers[15][0] ), .C1(n6171), .C2(
        \registers[14][0] ), .A(n5743), .ZN(n5742) );
  OAI22_X1 U1364 ( .A1(n2732), .A2(n6174), .B1(n4325), .B2(n6180), .ZN(n5743)
         );
  AOI221_X1 U1365 ( .B1(n6163), .B2(\registers[15][1] ), .C1(n6172), .C2(
        \registers[14][1] ), .A(n5711), .ZN(n5710) );
  OAI22_X1 U1366 ( .A1(n2733), .A2(n6175), .B1(n4326), .B2(n6181), .ZN(n5711)
         );
  AOI221_X1 U1367 ( .B1(n6166), .B2(\registers[15][3] ), .C1(n6170), .C2(
        \registers[14][3] ), .A(n5673), .ZN(n5672) );
  OAI22_X1 U1368 ( .A1(n2734), .A2(n6175), .B1(n4327), .B2(n6180), .ZN(n5673)
         );
  AOI221_X1 U1369 ( .B1(n6164), .B2(\registers[15][4] ), .C1(n6171), .C2(
        \registers[14][4] ), .A(n5654), .ZN(n5653) );
  OAI22_X1 U1370 ( .A1(n2735), .A2(n6176), .B1(n4328), .B2(n6181), .ZN(n5654)
         );
  AOI221_X1 U1371 ( .B1(n6165), .B2(\registers[15][6] ), .C1(n6172), .C2(
        \registers[14][6] ), .A(n5616), .ZN(n5615) );
  OAI22_X1 U1372 ( .A1(n2736), .A2(n6176), .B1(n4329), .B2(n6180), .ZN(n5616)
         );
  AOI221_X1 U1373 ( .B1(n6165), .B2(\registers[15][7] ), .C1(n6170), .C2(
        \registers[14][7] ), .A(n5597), .ZN(n5596) );
  OAI22_X1 U1374 ( .A1(n2737), .A2(n6177), .B1(n4330), .B2(n6181), .ZN(n5597)
         );
  AOI221_X1 U1375 ( .B1(n6167), .B2(\registers[15][9] ), .C1(n6171), .C2(
        \registers[14][9] ), .A(n5559), .ZN(n5558) );
  OAI22_X1 U1376 ( .A1(n2738), .A2(n6179), .B1(n4331), .B2(n6180), .ZN(n5559)
         );
  AOI221_X1 U1377 ( .B1(n6166), .B2(\registers[15][10] ), .C1(n6172), .C2(
        \registers[14][10] ), .A(n5540), .ZN(n5539) );
  OAI22_X1 U1378 ( .A1(n2739), .A2(n6174), .B1(n4332), .B2(n6181), .ZN(n5540)
         );
  AOI221_X1 U1379 ( .B1(n6168), .B2(\registers[15][12] ), .C1(n6170), .C2(
        \registers[14][12] ), .A(n5502), .ZN(n5501) );
  OAI22_X1 U1380 ( .A1(n2740), .A2(n6178), .B1(n4333), .B2(n6180), .ZN(n5502)
         );
  AOI221_X1 U1381 ( .B1(n6168), .B2(\registers[15][13] ), .C1(n6171), .C2(
        \registers[14][13] ), .A(n5483), .ZN(n5482) );
  OAI22_X1 U1382 ( .A1(n2741), .A2(n6179), .B1(n4334), .B2(n6181), .ZN(n5483)
         );
  AOI221_X1 U1383 ( .B1(n6167), .B2(\registers[15][15] ), .C1(n6172), .C2(
        \registers[14][15] ), .A(n5445), .ZN(n5444) );
  OAI22_X1 U1384 ( .A1(n2742), .A2(n6177), .B1(n4335), .B2(n6180), .ZN(n5445)
         );
  AOI221_X1 U1385 ( .B1(n6168), .B2(\registers[15][16] ), .C1(n6170), .C2(
        \registers[14][16] ), .A(n5426), .ZN(n5425) );
  OAI22_X1 U1386 ( .A1(n2743), .A2(n6178), .B1(n4336), .B2(n6181), .ZN(n5426)
         );
  AOI221_X1 U1387 ( .B1(n6169), .B2(\registers[15][18] ), .C1(n6171), .C2(
        \registers[14][18] ), .A(n5388), .ZN(n5387) );
  OAI22_X1 U1388 ( .A1(n2744), .A2(n6174), .B1(n4337), .B2(n6180), .ZN(n5388)
         );
  AOI221_X1 U1389 ( .B1(n6169), .B2(\registers[15][19] ), .C1(n6172), .C2(
        \registers[14][19] ), .A(n5369), .ZN(n5368) );
  OAI22_X1 U1390 ( .A1(n2745), .A2(n6175), .B1(n4338), .B2(n6181), .ZN(n5369)
         );
  AOI221_X1 U1391 ( .B1(n6169), .B2(\registers[15][21] ), .C1(n6170), .C2(
        \registers[14][21] ), .A(n5331), .ZN(n5330) );
  OAI22_X1 U1392 ( .A1(n2746), .A2(n6175), .B1(n4339), .B2(n6180), .ZN(n5331)
         );
  AOI221_X1 U1393 ( .B1(n6167), .B2(\registers[15][22] ), .C1(n6171), .C2(
        \registers[14][22] ), .A(n5312), .ZN(n5311) );
  OAI22_X1 U1394 ( .A1(n2747), .A2(n6176), .B1(n4340), .B2(n6181), .ZN(n5312)
         );
  AOI221_X1 U1395 ( .B1(n6163), .B2(\registers[15][24] ), .C1(n6172), .C2(
        \registers[14][24] ), .A(n5274), .ZN(n5273) );
  OAI22_X1 U1396 ( .A1(n2748), .A2(n6176), .B1(n4341), .B2(n6180), .ZN(n5274)
         );
  AOI221_X1 U1397 ( .B1(n6164), .B2(\registers[15][25] ), .C1(n6170), .C2(
        \registers[14][25] ), .A(n5255), .ZN(n5254) );
  OAI22_X1 U1398 ( .A1(n2749), .A2(n6177), .B1(n4342), .B2(n6181), .ZN(n5255)
         );
  AOI221_X1 U1399 ( .B1(n6164), .B2(\registers[15][27] ), .C1(n6171), .C2(
        \registers[14][27] ), .A(n5217), .ZN(n5216) );
  OAI22_X1 U1400 ( .A1(n2750), .A2(n6179), .B1(n4343), .B2(n6180), .ZN(n5217)
         );
  AOI221_X1 U1401 ( .B1(n6163), .B2(\registers[15][28] ), .C1(n6172), .C2(
        \registers[14][28] ), .A(n5198), .ZN(n5197) );
  OAI22_X1 U1402 ( .A1(n2751), .A2(n6174), .B1(n4344), .B2(n6181), .ZN(n5198)
         );
  AOI221_X1 U1403 ( .B1(n6165), .B2(\registers[15][30] ), .C1(n6170), .C2(
        \registers[14][30] ), .A(n5160), .ZN(n5159) );
  OAI22_X1 U1404 ( .A1(n2752), .A2(n6178), .B1(n4345), .B2(n6180), .ZN(n5160)
         );
  AOI221_X1 U1405 ( .B1(n6166), .B2(\registers[15][31] ), .C1(n6171), .C2(
        \registers[14][31] ), .A(n5127), .ZN(n5124) );
  OAI22_X1 U1406 ( .A1(n2753), .A2(n6179), .B1(n4346), .B2(n6181), .ZN(n5127)
         );
  AOI221_X1 U1407 ( .B1(n6372), .B2(\registers[15][0] ), .C1(n6380), .C2(
        \registers[14][0] ), .A(n5075), .ZN(n5074) );
  OAI22_X1 U1408 ( .A1(n2732), .A2(n6383), .B1(n4325), .B2(n6389), .ZN(n5075)
         );
  AOI221_X1 U1409 ( .B1(n6372), .B2(\registers[15][1] ), .C1(n6381), .C2(
        \registers[14][1] ), .A(n5042), .ZN(n5041) );
  OAI22_X1 U1410 ( .A1(n2733), .A2(n6384), .B1(n4326), .B2(n6390), .ZN(n5042)
         );
  AOI221_X1 U1411 ( .B1(n6374), .B2(\registers[15][3] ), .C1(n6379), .C2(
        \registers[14][3] ), .A(n5002), .ZN(n5001) );
  OAI22_X1 U1412 ( .A1(n2734), .A2(n6384), .B1(n4327), .B2(n6389), .ZN(n5002)
         );
  AOI221_X1 U1413 ( .B1(n6374), .B2(\registers[15][4] ), .C1(n6380), .C2(
        \registers[14][4] ), .A(n4982), .ZN(n4981) );
  OAI22_X1 U1414 ( .A1(n2735), .A2(n6385), .B1(n4328), .B2(n6390), .ZN(n4982)
         );
  AOI221_X1 U1415 ( .B1(n6375), .B2(\registers[15][6] ), .C1(n6381), .C2(
        \registers[14][6] ), .A(n4942), .ZN(n4941) );
  OAI22_X1 U1416 ( .A1(n2736), .A2(n6385), .B1(n4329), .B2(n6389), .ZN(n4942)
         );
  AOI221_X1 U1417 ( .B1(n6376), .B2(\registers[15][7] ), .C1(n6379), .C2(
        \registers[14][7] ), .A(n4922), .ZN(n4921) );
  OAI22_X1 U1418 ( .A1(n2737), .A2(n6386), .B1(n4330), .B2(n6390), .ZN(n4922)
         );
  AOI221_X1 U1419 ( .B1(n6376), .B2(\registers[15][9] ), .C1(n6380), .C2(
        \registers[14][9] ), .A(n4882), .ZN(n4881) );
  OAI22_X1 U1420 ( .A1(n2738), .A2(n6388), .B1(n4331), .B2(n6389), .ZN(n4882)
         );
  AOI221_X1 U1421 ( .B1(n6376), .B2(\registers[15][10] ), .C1(n6381), .C2(
        \registers[14][10] ), .A(n4862), .ZN(n4861) );
  OAI22_X1 U1422 ( .A1(n2739), .A2(n6383), .B1(n4332), .B2(n6390), .ZN(n4862)
         );
  AOI221_X1 U1423 ( .B1(n6377), .B2(\registers[15][12] ), .C1(n6379), .C2(
        \registers[14][12] ), .A(n4822), .ZN(n4821) );
  OAI22_X1 U1424 ( .A1(n2740), .A2(n6387), .B1(n4333), .B2(n6389), .ZN(n4822)
         );
  AOI221_X1 U1425 ( .B1(n6377), .B2(\registers[15][13] ), .C1(n6380), .C2(
        \registers[14][13] ), .A(n4802), .ZN(n4801) );
  OAI22_X1 U1426 ( .A1(n2741), .A2(n6388), .B1(n4334), .B2(n6390), .ZN(n4802)
         );
  AOI221_X1 U1427 ( .B1(n6376), .B2(\registers[15][15] ), .C1(n6381), .C2(
        \registers[14][15] ), .A(n4762), .ZN(n4761) );
  OAI22_X1 U1428 ( .A1(n2742), .A2(n6386), .B1(n4335), .B2(n6389), .ZN(n4762)
         );
  AOI221_X1 U1429 ( .B1(n6377), .B2(\registers[15][16] ), .C1(n6379), .C2(
        \registers[14][16] ), .A(n4742), .ZN(n4741) );
  OAI22_X1 U1430 ( .A1(n2743), .A2(n6387), .B1(n4336), .B2(n6390), .ZN(n4742)
         );
  AOI221_X1 U1431 ( .B1(n6378), .B2(\registers[15][18] ), .C1(n6380), .C2(
        \registers[14][18] ), .A(n4702), .ZN(n4701) );
  OAI22_X1 U1432 ( .A1(n2744), .A2(n6383), .B1(n4337), .B2(n6389), .ZN(n4702)
         );
  AOI221_X1 U1433 ( .B1(n6378), .B2(\registers[15][19] ), .C1(n6381), .C2(
        \registers[14][19] ), .A(n4682), .ZN(n4681) );
  OAI22_X1 U1434 ( .A1(n2745), .A2(n6384), .B1(n4338), .B2(n6390), .ZN(n4682)
         );
  AOI221_X1 U1435 ( .B1(n6378), .B2(\registers[15][21] ), .C1(n6379), .C2(
        \registers[14][21] ), .A(n4642), .ZN(n4641) );
  OAI22_X1 U1436 ( .A1(n2746), .A2(n6384), .B1(n4339), .B2(n6389), .ZN(n4642)
         );
  AOI221_X1 U1437 ( .B1(n6372), .B2(\registers[15][22] ), .C1(n6380), .C2(
        \registers[14][22] ), .A(n4622), .ZN(n4621) );
  OAI22_X1 U1438 ( .A1(n2747), .A2(n6385), .B1(n4340), .B2(n6390), .ZN(n4622)
         );
  AOI221_X1 U1439 ( .B1(n6373), .B2(\registers[15][24] ), .C1(n6381), .C2(
        \registers[14][24] ), .A(n4582), .ZN(n4581) );
  OAI22_X1 U1440 ( .A1(n2748), .A2(n6385), .B1(n4341), .B2(n6389), .ZN(n4582)
         );
  AOI221_X1 U1441 ( .B1(n6374), .B2(\registers[15][25] ), .C1(n6379), .C2(
        \registers[14][25] ), .A(n4562), .ZN(n4561) );
  OAI22_X1 U1442 ( .A1(n2749), .A2(n6386), .B1(n4342), .B2(n6390), .ZN(n4562)
         );
  AOI221_X1 U1443 ( .B1(n6375), .B2(\registers[15][27] ), .C1(n6380), .C2(
        \registers[14][27] ), .A(n4522), .ZN(n4521) );
  OAI22_X1 U1444 ( .A1(n2750), .A2(n6388), .B1(n4343), .B2(n6389), .ZN(n4522)
         );
  AOI221_X1 U1445 ( .B1(n6375), .B2(\registers[15][28] ), .C1(n6381), .C2(
        \registers[14][28] ), .A(n4502), .ZN(n4501) );
  OAI22_X1 U1446 ( .A1(n2751), .A2(n6383), .B1(n4344), .B2(n6390), .ZN(n4502)
         );
  AOI221_X1 U1447 ( .B1(n6378), .B2(\registers[15][30] ), .C1(n6379), .C2(
        \registers[14][30] ), .A(n4462), .ZN(n4461) );
  OAI22_X1 U1448 ( .A1(n2752), .A2(n6387), .B1(n4345), .B2(n6389), .ZN(n4462)
         );
  AOI221_X1 U1449 ( .B1(n6376), .B2(\registers[15][31] ), .C1(n6380), .C2(
        \registers[14][31] ), .A(n4428), .ZN(n4425) );
  OAI22_X1 U1450 ( .A1(n2753), .A2(n6388), .B1(n4346), .B2(n6390), .ZN(n4428)
         );
  AOI221_X1 U1451 ( .B1(n6262), .B2(\registers[5][4] ), .C1(n6264), .C2(
        \registers[4][4] ), .A(n5646), .ZN(n5645) );
  OAI22_X1 U1452 ( .A1(n2754), .A2(n6268), .B1(n4347), .B2(n6273), .ZN(n5646)
         );
  AOI221_X1 U1453 ( .B1(n6261), .B2(\registers[5][6] ), .C1(n6263), .C2(
        \registers[4][6] ), .A(n5608), .ZN(n5607) );
  OAI22_X1 U1454 ( .A1(n2758), .A2(n6268), .B1(n4348), .B2(n6272), .ZN(n5608)
         );
  AOI221_X1 U1455 ( .B1(n6262), .B2(\registers[5][7] ), .C1(n6264), .C2(
        \registers[4][7] ), .A(n5589), .ZN(n5588) );
  OAI22_X1 U1456 ( .A1(n2759), .A2(n6269), .B1(n4349), .B2(n6273), .ZN(n5589)
         );
  AOI221_X1 U1457 ( .B1(n6261), .B2(\registers[5][9] ), .C1(n6263), .C2(
        \registers[4][9] ), .A(n5551), .ZN(n5550) );
  OAI22_X1 U1458 ( .A1(n2760), .A2(n6271), .B1(n4350), .B2(n6272), .ZN(n5551)
         );
  AOI221_X1 U1459 ( .B1(n6261), .B2(\registers[5][12] ), .C1(n6263), .C2(
        \registers[4][12] ), .A(n5494), .ZN(n5493) );
  OAI22_X1 U1460 ( .A1(n2761), .A2(n6270), .B1(n4351), .B2(n6272), .ZN(n5494)
         );
  AOI221_X1 U1461 ( .B1(n6262), .B2(\registers[5][13] ), .C1(n6264), .C2(
        \registers[4][13] ), .A(n5475), .ZN(n5474) );
  OAI22_X1 U1462 ( .A1(n2762), .A2(n6271), .B1(n4352), .B2(n6273), .ZN(n5475)
         );
  AOI221_X1 U1463 ( .B1(n6261), .B2(\registers[5][15] ), .C1(n6263), .C2(
        \registers[4][15] ), .A(n5437), .ZN(n5436) );
  OAI22_X1 U1464 ( .A1(n2763), .A2(n6269), .B1(n4353), .B2(n6272), .ZN(n5437)
         );
  AOI221_X1 U1465 ( .B1(n6262), .B2(\registers[5][16] ), .C1(n6264), .C2(
        \registers[4][16] ), .A(n5418), .ZN(n5417) );
  OAI22_X1 U1466 ( .A1(n2764), .A2(n6270), .B1(n4356), .B2(n6273), .ZN(n5418)
         );
  AOI221_X1 U1467 ( .B1(n6262), .B2(\registers[5][22] ), .C1(n6264), .C2(
        \registers[4][22] ), .A(n5304), .ZN(n5303) );
  OAI22_X1 U1468 ( .A1(n2765), .A2(n6268), .B1(n4390), .B2(n6273), .ZN(n5304)
         );
  AOI221_X1 U1469 ( .B1(n6261), .B2(\registers[5][24] ), .C1(n6263), .C2(
        \registers[4][24] ), .A(n5266), .ZN(n5265) );
  OAI22_X1 U1470 ( .A1(n2766), .A2(n6268), .B1(n5759), .B2(n6272), .ZN(n5266)
         );
  AOI221_X1 U1471 ( .B1(n6262), .B2(\registers[5][25] ), .C1(n6264), .C2(
        \registers[4][25] ), .A(n5247), .ZN(n5246) );
  OAI22_X1 U1472 ( .A1(n2767), .A2(n6269), .B1(n5760), .B2(n6273), .ZN(n5247)
         );
  AOI221_X1 U1473 ( .B1(n6261), .B2(\registers[5][27] ), .C1(n6263), .C2(
        \registers[4][27] ), .A(n5209), .ZN(n5208) );
  OAI22_X1 U1474 ( .A1(n2768), .A2(n6271), .B1(n5761), .B2(n6272), .ZN(n5209)
         );
  AOI221_X1 U1475 ( .B1(n6261), .B2(\registers[5][30] ), .C1(n6263), .C2(
        \registers[4][30] ), .A(n5152), .ZN(n5151) );
  OAI22_X1 U1476 ( .A1(n2769), .A2(n6270), .B1(n5762), .B2(n6272), .ZN(n5152)
         );
  AOI221_X1 U1477 ( .B1(n6262), .B2(\registers[5][31] ), .C1(n6264), .C2(
        \registers[4][31] ), .A(n5103), .ZN(n5100) );
  OAI22_X1 U1478 ( .A1(n2770), .A2(n6271), .B1(n5763), .B2(n6273), .ZN(n5103)
         );
  AOI221_X1 U1479 ( .B1(n6373), .B2(\registers[15][2] ), .C1(n6379), .C2(
        \registers[14][2] ), .A(n5022), .ZN(n5021) );
  OAI22_X1 U1480 ( .A1(n2771), .A2(n6383), .B1(n5764), .B2(n4430), .ZN(n5022)
         );
  AOI221_X1 U1481 ( .B1(n6374), .B2(\registers[15][5] ), .C1(n6380), .C2(
        \registers[14][5] ), .A(n4962), .ZN(n4961) );
  OAI22_X1 U1482 ( .A1(n2772), .A2(n6386), .B1(n5765), .B2(n4430), .ZN(n4962)
         );
  AOI221_X1 U1483 ( .B1(n6374), .B2(\registers[15][8] ), .C1(n6381), .C2(
        \registers[14][8] ), .A(n4902), .ZN(n4901) );
  OAI22_X1 U1484 ( .A1(n2773), .A2(n6387), .B1(n5766), .B2(n4430), .ZN(n4902)
         );
  AOI221_X1 U1485 ( .B1(n6373), .B2(\registers[15][11] ), .C1(n6379), .C2(
        \registers[14][11] ), .A(n4842), .ZN(n4841) );
  OAI22_X1 U1486 ( .A1(n2774), .A2(n6384), .B1(n5767), .B2(n4430), .ZN(n4842)
         );
  AOI221_X1 U1487 ( .B1(n6373), .B2(\registers[15][14] ), .C1(n6380), .C2(
        \registers[14][14] ), .A(n4782), .ZN(n4781) );
  OAI22_X1 U1488 ( .A1(n2775), .A2(n6385), .B1(n5768), .B2(n4430), .ZN(n4782)
         );
  AOI221_X1 U1489 ( .B1(n6377), .B2(\registers[15][17] ), .C1(n6381), .C2(
        \registers[14][17] ), .A(n4722), .ZN(n4721) );
  OAI22_X1 U1490 ( .A1(n2776), .A2(n6388), .B1(n5769), .B2(n4430), .ZN(n4722)
         );
  AOI221_X1 U1491 ( .B1(n6378), .B2(\registers[15][20] ), .C1(n6379), .C2(
        \registers[14][20] ), .A(n4662), .ZN(n4661) );
  OAI22_X1 U1492 ( .A1(n2777), .A2(n6383), .B1(n5770), .B2(n4430), .ZN(n4662)
         );
  AOI221_X1 U1493 ( .B1(n6373), .B2(\registers[15][23] ), .C1(n6380), .C2(
        \registers[14][23] ), .A(n4602), .ZN(n4601) );
  OAI22_X1 U1494 ( .A1(n2778), .A2(n6386), .B1(n5771), .B2(n4430), .ZN(n4602)
         );
  AOI221_X1 U1495 ( .B1(n6372), .B2(\registers[15][26] ), .C1(n6381), .C2(
        \registers[14][26] ), .A(n4542), .ZN(n4541) );
  OAI22_X1 U1496 ( .A1(n2779), .A2(n6387), .B1(n5772), .B2(n4430), .ZN(n4542)
         );
  AOI221_X1 U1497 ( .B1(n6375), .B2(\registers[15][29] ), .C1(n6379), .C2(
        \registers[14][29] ), .A(n4482), .ZN(n4481) );
  OAI22_X1 U1498 ( .A1(n2780), .A2(n6384), .B1(n5773), .B2(n4430), .ZN(n4482)
         );
  AOI221_X1 U1499 ( .B1(n5101), .B2(\registers[5][2] ), .C1(n5102), .C2(
        \registers[4][2] ), .A(n5684), .ZN(n5683) );
  OAI22_X1 U1500 ( .A1(n2781), .A2(n6266), .B1(n5774), .B2(n5105), .ZN(n5684)
         );
  AOI221_X1 U1501 ( .B1(n5101), .B2(\registers[5][5] ), .C1(n5102), .C2(
        \registers[4][5] ), .A(n5627), .ZN(n5626) );
  OAI22_X1 U1502 ( .A1(n2782), .A2(n6269), .B1(n5775), .B2(n5105), .ZN(n5627)
         );
  AOI221_X1 U1503 ( .B1(n5101), .B2(\registers[5][8] ), .C1(n5102), .C2(
        \registers[4][8] ), .A(n5570), .ZN(n5569) );
  OAI22_X1 U1504 ( .A1(n2783), .A2(n6270), .B1(n5776), .B2(n5105), .ZN(n5570)
         );
  AOI221_X1 U1505 ( .B1(n5101), .B2(\registers[5][11] ), .C1(n5102), .C2(
        \registers[4][11] ), .A(n5513), .ZN(n5512) );
  OAI22_X1 U1506 ( .A1(n2784), .A2(n6267), .B1(n5777), .B2(n5105), .ZN(n5513)
         );
  AOI221_X1 U1507 ( .B1(n5101), .B2(\registers[5][14] ), .C1(n5102), .C2(
        \registers[4][14] ), .A(n5456), .ZN(n5455) );
  OAI22_X1 U1508 ( .A1(n2785), .A2(n6268), .B1(n5778), .B2(n5105), .ZN(n5456)
         );
  AOI221_X1 U1509 ( .B1(n5101), .B2(\registers[5][17] ), .C1(n5102), .C2(
        \registers[4][17] ), .A(n5399), .ZN(n5398) );
  OAI22_X1 U1510 ( .A1(n2786), .A2(n6271), .B1(n5779), .B2(n5105), .ZN(n5399)
         );
  AOI221_X1 U1511 ( .B1(n5101), .B2(\registers[5][20] ), .C1(n5102), .C2(
        \registers[4][20] ), .A(n5342), .ZN(n5341) );
  OAI22_X1 U1512 ( .A1(n2787), .A2(n6266), .B1(n5780), .B2(n5105), .ZN(n5342)
         );
  AOI221_X1 U1513 ( .B1(n5101), .B2(\registers[5][23] ), .C1(n5102), .C2(
        \registers[4][23] ), .A(n5285), .ZN(n5284) );
  OAI22_X1 U1514 ( .A1(n2788), .A2(n6269), .B1(n5781), .B2(n5105), .ZN(n5285)
         );
  AOI221_X1 U1515 ( .B1(n5101), .B2(\registers[5][26] ), .C1(n5102), .C2(
        \registers[4][26] ), .A(n5228), .ZN(n5227) );
  OAI22_X1 U1516 ( .A1(n2789), .A2(n6270), .B1(n5782), .B2(n5105), .ZN(n5228)
         );
  AOI221_X1 U1517 ( .B1(n5101), .B2(\registers[5][29] ), .C1(n5102), .C2(
        \registers[4][29] ), .A(n5171), .ZN(n5170) );
  OAI22_X1 U1518 ( .A1(n2791), .A2(n6267), .B1(n5783), .B2(n5105), .ZN(n5171)
         );
  AOI221_X1 U1519 ( .B1(n6412), .B2(\registers[21][0] ), .C1(n6420), .C2(
        \registers[20][0] ), .A(n5063), .ZN(n5052) );
  OAI22_X1 U1520 ( .A1(n2793), .A2(n6423), .B1(n5785), .B2(n6429), .ZN(n5063)
         );
  AOI221_X1 U1521 ( .B1(n6413), .B2(\registers[21][1] ), .C1(n6421), .C2(
        \registers[20][1] ), .A(n5036), .ZN(n5031) );
  OAI22_X1 U1522 ( .A1(n2795), .A2(n6424), .B1(n5787), .B2(n6430), .ZN(n5036)
         );
  AOI221_X1 U1523 ( .B1(n6414), .B2(\registers[21][3] ), .C1(n6419), .C2(
        \registers[20][3] ), .A(n4996), .ZN(n4991) );
  OAI22_X1 U1524 ( .A1(n2799), .A2(n6424), .B1(n5791), .B2(n6429), .ZN(n4996)
         );
  AOI221_X1 U1525 ( .B1(n6414), .B2(\registers[21][4] ), .C1(n6420), .C2(
        \registers[20][4] ), .A(n4976), .ZN(n4971) );
  OAI22_X1 U1526 ( .A1(n2801), .A2(n6425), .B1(n5793), .B2(n6430), .ZN(n4976)
         );
  AOI221_X1 U1527 ( .B1(n6415), .B2(\registers[21][6] ), .C1(n6421), .C2(
        \registers[20][6] ), .A(n4936), .ZN(n4931) );
  OAI22_X1 U1528 ( .A1(n2805), .A2(n6425), .B1(n5797), .B2(n6429), .ZN(n4936)
         );
  AOI221_X1 U1529 ( .B1(n6418), .B2(\registers[21][7] ), .C1(n6419), .C2(
        \registers[20][7] ), .A(n4916), .ZN(n4911) );
  OAI22_X1 U1530 ( .A1(n2807), .A2(n6426), .B1(n5799), .B2(n6430), .ZN(n4916)
         );
  AOI221_X1 U1531 ( .B1(n6416), .B2(\registers[21][9] ), .C1(n6420), .C2(
        \registers[20][9] ), .A(n4876), .ZN(n4871) );
  OAI22_X1 U1532 ( .A1(n2811), .A2(n6428), .B1(n5803), .B2(n6429), .ZN(n4876)
         );
  AOI221_X1 U1533 ( .B1(n6416), .B2(\registers[21][10] ), .C1(n6421), .C2(
        \registers[20][10] ), .A(n4856), .ZN(n4851) );
  OAI22_X1 U1534 ( .A1(n2813), .A2(n6423), .B1(n5805), .B2(n6430), .ZN(n4856)
         );
  AOI221_X1 U1535 ( .B1(n6417), .B2(\registers[21][12] ), .C1(n6419), .C2(
        \registers[20][12] ), .A(n4816), .ZN(n4811) );
  OAI22_X1 U1536 ( .A1(n2817), .A2(n6427), .B1(n5809), .B2(n6429), .ZN(n4816)
         );
  AOI221_X1 U1537 ( .B1(n6417), .B2(\registers[21][13] ), .C1(n6420), .C2(
        \registers[20][13] ), .A(n4796), .ZN(n4791) );
  OAI22_X1 U1538 ( .A1(n2819), .A2(n6428), .B1(n5811), .B2(n6430), .ZN(n4796)
         );
  AOI221_X1 U1539 ( .B1(n6413), .B2(\registers[21][15] ), .C1(n6421), .C2(
        \registers[20][15] ), .A(n4756), .ZN(n4751) );
  OAI22_X1 U1540 ( .A1(n2823), .A2(n6426), .B1(n5815), .B2(n6429), .ZN(n4756)
         );
  AOI221_X1 U1541 ( .B1(n6417), .B2(\registers[21][16] ), .C1(n6419), .C2(
        \registers[20][16] ), .A(n4736), .ZN(n4731) );
  OAI22_X1 U1542 ( .A1(n2827), .A2(n6427), .B1(n5817), .B2(n6430), .ZN(n4736)
         );
  AOI221_X1 U1543 ( .B1(n6418), .B2(\registers[21][18] ), .C1(n6420), .C2(
        \registers[20][18] ), .A(n4696), .ZN(n4691) );
  OAI22_X1 U1544 ( .A1(n2831), .A2(n6423), .B1(n5821), .B2(n6429), .ZN(n4696)
         );
  AOI221_X1 U1545 ( .B1(n6418), .B2(\registers[21][19] ), .C1(n6421), .C2(
        \registers[20][19] ), .A(n4676), .ZN(n4671) );
  OAI22_X1 U1546 ( .A1(n2833), .A2(n6424), .B1(n5823), .B2(n6430), .ZN(n4676)
         );
  AOI221_X1 U1547 ( .B1(n6418), .B2(\registers[21][21] ), .C1(n6419), .C2(
        \registers[20][21] ), .A(n4636), .ZN(n4631) );
  OAI22_X1 U1548 ( .A1(n2837), .A2(n6424), .B1(n5827), .B2(n6429), .ZN(n4636)
         );
  AOI221_X1 U1549 ( .B1(n6412), .B2(\registers[21][22] ), .C1(n6420), .C2(
        \registers[20][22] ), .A(n4616), .ZN(n4611) );
  OAI22_X1 U1550 ( .A1(n4213), .A2(n6425), .B1(n5912), .B2(n6430), .ZN(n4616)
         );
  AOI221_X1 U1551 ( .B1(n6413), .B2(\registers[21][24] ), .C1(n6421), .C2(
        \registers[20][24] ), .A(n4576), .ZN(n4571) );
  OAI22_X1 U1552 ( .A1(n4215), .A2(n6425), .B1(n5914), .B2(n6429), .ZN(n4576)
         );
  AOI221_X1 U1553 ( .B1(n6414), .B2(\registers[21][25] ), .C1(n6419), .C2(
        \registers[20][25] ), .A(n4556), .ZN(n4551) );
  OAI22_X1 U1554 ( .A1(n4216), .A2(n6426), .B1(n5915), .B2(n6430), .ZN(n4556)
         );
  AOI221_X1 U1555 ( .B1(n6414), .B2(\registers[21][27] ), .C1(n6420), .C2(
        \registers[20][27] ), .A(n4516), .ZN(n4511) );
  OAI22_X1 U1556 ( .A1(n4219), .A2(n6428), .B1(n5917), .B2(n6429), .ZN(n4516)
         );
  AOI221_X1 U1557 ( .B1(n6415), .B2(\registers[21][28] ), .C1(n6421), .C2(
        \registers[20][28] ), .A(n4496), .ZN(n4491) );
  OAI22_X1 U1558 ( .A1(n2845), .A2(n6423), .B1(n5835), .B2(n6430), .ZN(n4496)
         );
  AOI221_X1 U1559 ( .B1(n6416), .B2(\registers[21][30] ), .C1(n6419), .C2(
        \registers[20][30] ), .A(n4456), .ZN(n4451) );
  OAI22_X1 U1560 ( .A1(n2849), .A2(n6427), .B1(n5839), .B2(n6429), .ZN(n4456)
         );
  AOI221_X1 U1561 ( .B1(n6416), .B2(\registers[21][31] ), .C1(n6420), .C2(
        \registers[20][31] ), .A(n4414), .ZN(n4399) );
  OAI22_X1 U1562 ( .A1(n2851), .A2(n6428), .B1(n5841), .B2(n6430), .ZN(n4414)
         );
  AOI221_X1 U1563 ( .B1(n6413), .B2(\registers[21][2] ), .C1(n6419), .C2(
        \registers[20][2] ), .A(n5016), .ZN(n5011) );
  OAI22_X1 U1564 ( .A1(n2797), .A2(n6423), .B1(n5789), .B2(n4416), .ZN(n5016)
         );
  AOI221_X1 U1565 ( .B1(n6412), .B2(\registers[21][5] ), .C1(n6420), .C2(
        \registers[20][5] ), .A(n4956), .ZN(n4951) );
  OAI22_X1 U1566 ( .A1(n2803), .A2(n6426), .B1(n5795), .B2(n4416), .ZN(n4956)
         );
  AOI221_X1 U1567 ( .B1(n6415), .B2(\registers[21][8] ), .C1(n6421), .C2(
        \registers[20][8] ), .A(n4896), .ZN(n4891) );
  OAI22_X1 U1568 ( .A1(n2809), .A2(n6427), .B1(n5801), .B2(n4416), .ZN(n4896)
         );
  AOI221_X1 U1569 ( .B1(n6413), .B2(\registers[21][11] ), .C1(n6419), .C2(
        \registers[20][11] ), .A(n4836), .ZN(n4831) );
  OAI22_X1 U1570 ( .A1(n2815), .A2(n6424), .B1(n5807), .B2(n4416), .ZN(n4836)
         );
  AOI221_X1 U1571 ( .B1(n6416), .B2(\registers[21][14] ), .C1(n6420), .C2(
        \registers[20][14] ), .A(n4776), .ZN(n4771) );
  OAI22_X1 U1572 ( .A1(n2821), .A2(n6425), .B1(n5813), .B2(n4416), .ZN(n4776)
         );
  AOI221_X1 U1573 ( .B1(n6417), .B2(\registers[21][17] ), .C1(n6421), .C2(
        \registers[20][17] ), .A(n4716), .ZN(n4711) );
  OAI22_X1 U1574 ( .A1(n2829), .A2(n6428), .B1(n5819), .B2(n4416), .ZN(n4716)
         );
  AOI221_X1 U1575 ( .B1(n6418), .B2(\registers[21][20] ), .C1(n6419), .C2(
        \registers[20][20] ), .A(n4656), .ZN(n4651) );
  OAI22_X1 U1576 ( .A1(n2835), .A2(n6423), .B1(n5825), .B2(n4416), .ZN(n4656)
         );
  AOI221_X1 U1577 ( .B1(n6412), .B2(\registers[21][23] ), .C1(n6420), .C2(
        \registers[20][23] ), .A(n4596), .ZN(n4591) );
  OAI22_X1 U1578 ( .A1(n4214), .A2(n6426), .B1(n5913), .B2(n4416), .ZN(n4596)
         );
  AOI221_X1 U1579 ( .B1(n6415), .B2(\registers[21][26] ), .C1(n6421), .C2(
        \registers[20][26] ), .A(n4536), .ZN(n4531) );
  OAI22_X1 U1580 ( .A1(n4218), .A2(n6427), .B1(n5916), .B2(n4416), .ZN(n4536)
         );
  AOI221_X1 U1581 ( .B1(n6415), .B2(\registers[21][29] ), .C1(n6419), .C2(
        \registers[20][29] ), .A(n4476), .ZN(n4471) );
  OAI22_X1 U1582 ( .A1(n2847), .A2(n6424), .B1(n5837), .B2(n4416), .ZN(n4476)
         );
  OAI221_X1 U1583 ( .B1(n6073), .B2(n3050), .C1(n1748), .C2(n6074), .A(n5715), 
        .ZN(n3051) );
  OAI21_X1 U1584 ( .B1(n5716), .B2(n5717), .A(n6275), .ZN(n5715) );
  NAND4_X1 U1585 ( .A1(n5739), .A2(n5740), .A3(n5741), .A4(n5742), .ZN(n5716)
         );
  NAND4_X1 U1586 ( .A1(n5719), .A2(n5720), .A3(n5721), .A4(n5722), .ZN(n5717)
         );
  OAI221_X1 U1587 ( .B1(n5091), .B2(n3049), .C1(n1746), .C2(n6075), .A(n5696), 
        .ZN(n3052) );
  OAI21_X1 U1588 ( .B1(n5697), .B2(n5698), .A(n6276), .ZN(n5696) );
  NAND4_X1 U1589 ( .A1(n5707), .A2(n5708), .A3(n5709), .A4(n5710), .ZN(n5697)
         );
  NAND4_X1 U1590 ( .A1(n5699), .A2(n5700), .A3(n5701), .A4(n5702), .ZN(n5698)
         );
  OAI221_X1 U1591 ( .B1(n6073), .B2(n3047), .C1(n1742), .C2(n6074), .A(n5658), 
        .ZN(n3054) );
  OAI21_X1 U1592 ( .B1(n5659), .B2(n5660), .A(n6274), .ZN(n5658) );
  NAND4_X1 U1593 ( .A1(n5669), .A2(n5670), .A3(n5671), .A4(n5672), .ZN(n5659)
         );
  NAND4_X1 U1594 ( .A1(n5661), .A2(n5662), .A3(n5663), .A4(n5664), .ZN(n5660)
         );
  OAI221_X1 U1595 ( .B1(n5091), .B2(n3046), .C1(n1740), .C2(n6075), .A(n5639), 
        .ZN(n3055) );
  OAI21_X1 U1596 ( .B1(n5640), .B2(n5641), .A(n6275), .ZN(n5639) );
  NAND4_X1 U1597 ( .A1(n5650), .A2(n5651), .A3(n5652), .A4(n5653), .ZN(n5640)
         );
  NAND4_X1 U1598 ( .A1(n5642), .A2(n5643), .A3(n5644), .A4(n5645), .ZN(n5641)
         );
  OAI221_X1 U1599 ( .B1(n6073), .B2(n3044), .C1(n1736), .C2(n6074), .A(n5601), 
        .ZN(n3057) );
  OAI21_X1 U1600 ( .B1(n5602), .B2(n5603), .A(n6276), .ZN(n5601) );
  NAND4_X1 U1601 ( .A1(n5612), .A2(n5613), .A3(n5614), .A4(n5615), .ZN(n5602)
         );
  NAND4_X1 U1602 ( .A1(n5604), .A2(n5605), .A3(n5606), .A4(n5607), .ZN(n5603)
         );
  OAI221_X1 U1603 ( .B1(n5091), .B2(n3043), .C1(n1734), .C2(n6075), .A(n5582), 
        .ZN(n3058) );
  OAI21_X1 U1604 ( .B1(n5583), .B2(n5584), .A(n6274), .ZN(n5582) );
  NAND4_X1 U1605 ( .A1(n5593), .A2(n5594), .A3(n5595), .A4(n5596), .ZN(n5583)
         );
  NAND4_X1 U1606 ( .A1(n5585), .A2(n5586), .A3(n5587), .A4(n5588), .ZN(n5584)
         );
  OAI221_X1 U1607 ( .B1(n6073), .B2(n3041), .C1(n1730), .C2(n6074), .A(n5544), 
        .ZN(n3060) );
  OAI21_X1 U1608 ( .B1(n5545), .B2(n5546), .A(n6275), .ZN(n5544) );
  NAND4_X1 U1609 ( .A1(n5555), .A2(n5556), .A3(n5557), .A4(n5558), .ZN(n5545)
         );
  NAND4_X1 U1610 ( .A1(n5547), .A2(n5548), .A3(n5549), .A4(n5550), .ZN(n5546)
         );
  OAI221_X1 U1611 ( .B1(n5091), .B2(n3040), .C1(n1728), .C2(n6075), .A(n5525), 
        .ZN(n3061) );
  OAI21_X1 U1612 ( .B1(n5526), .B2(n5527), .A(n6276), .ZN(n5525) );
  NAND4_X1 U1613 ( .A1(n5536), .A2(n5537), .A3(n5538), .A4(n5539), .ZN(n5526)
         );
  NAND4_X1 U1614 ( .A1(n5528), .A2(n5529), .A3(n5530), .A4(n5531), .ZN(n5527)
         );
  OAI221_X1 U1615 ( .B1(n6073), .B2(n3038), .C1(n1724), .C2(n6074), .A(n5487), 
        .ZN(n3063) );
  OAI21_X1 U1616 ( .B1(n5488), .B2(n5489), .A(n6274), .ZN(n5487) );
  NAND4_X1 U1617 ( .A1(n5498), .A2(n5499), .A3(n5500), .A4(n5501), .ZN(n5488)
         );
  NAND4_X1 U1618 ( .A1(n5490), .A2(n5491), .A3(n5492), .A4(n5493), .ZN(n5489)
         );
  OAI221_X1 U1619 ( .B1(n5091), .B2(n3037), .C1(n1722), .C2(n6075), .A(n5468), 
        .ZN(n3064) );
  OAI21_X1 U1620 ( .B1(n5469), .B2(n5470), .A(n6275), .ZN(n5468) );
  NAND4_X1 U1621 ( .A1(n5479), .A2(n5480), .A3(n5481), .A4(n5482), .ZN(n5469)
         );
  NAND4_X1 U1622 ( .A1(n5471), .A2(n5472), .A3(n5473), .A4(n5474), .ZN(n5470)
         );
  OAI221_X1 U1623 ( .B1(n6073), .B2(n3035), .C1(n1718), .C2(n6074), .A(n5430), 
        .ZN(n3066) );
  OAI21_X1 U1624 ( .B1(n5431), .B2(n5432), .A(n6276), .ZN(n5430) );
  NAND4_X1 U1625 ( .A1(n5441), .A2(n5442), .A3(n5443), .A4(n5444), .ZN(n5431)
         );
  NAND4_X1 U1626 ( .A1(n5433), .A2(n5434), .A3(n5435), .A4(n5436), .ZN(n5432)
         );
  OAI221_X1 U1627 ( .B1(n5091), .B2(n3034), .C1(n1716), .C2(n6075), .A(n5411), 
        .ZN(n3067) );
  OAI21_X1 U1628 ( .B1(n5412), .B2(n5413), .A(n6274), .ZN(n5411) );
  NAND4_X1 U1629 ( .A1(n5422), .A2(n5423), .A3(n5424), .A4(n5425), .ZN(n5412)
         );
  NAND4_X1 U1630 ( .A1(n5414), .A2(n5415), .A3(n5416), .A4(n5417), .ZN(n5413)
         );
  OAI221_X1 U1631 ( .B1(n6073), .B2(n3032), .C1(n1712), .C2(n6074), .A(n5373), 
        .ZN(n3069) );
  OAI21_X1 U1632 ( .B1(n5374), .B2(n5375), .A(n6275), .ZN(n5373) );
  NAND4_X1 U1633 ( .A1(n5384), .A2(n5385), .A3(n5386), .A4(n5387), .ZN(n5374)
         );
  NAND4_X1 U1634 ( .A1(n5376), .A2(n5377), .A3(n5378), .A4(n5379), .ZN(n5375)
         );
  OAI221_X1 U1635 ( .B1(n5091), .B2(n3031), .C1(n1710), .C2(n6075), .A(n5354), 
        .ZN(n3070) );
  OAI21_X1 U1636 ( .B1(n5355), .B2(n5356), .A(n6276), .ZN(n5354) );
  NAND4_X1 U1637 ( .A1(n5365), .A2(n5366), .A3(n5367), .A4(n5368), .ZN(n5355)
         );
  NAND4_X1 U1638 ( .A1(n5357), .A2(n5358), .A3(n5359), .A4(n5360), .ZN(n5356)
         );
  OAI221_X1 U1639 ( .B1(n6073), .B2(n3029), .C1(n1706), .C2(n6074), .A(n5316), 
        .ZN(n3072) );
  OAI21_X1 U1640 ( .B1(n5317), .B2(n5318), .A(n6274), .ZN(n5316) );
  NAND4_X1 U1641 ( .A1(n5327), .A2(n5328), .A3(n5329), .A4(n5330), .ZN(n5317)
         );
  NAND4_X1 U1642 ( .A1(n5319), .A2(n5320), .A3(n5321), .A4(n5322), .ZN(n5318)
         );
  OAI221_X1 U1643 ( .B1(n5091), .B2(n3028), .C1(n1704), .C2(n6075), .A(n5297), 
        .ZN(n3073) );
  OAI21_X1 U1644 ( .B1(n5298), .B2(n5299), .A(n6275), .ZN(n5297) );
  NAND4_X1 U1645 ( .A1(n5308), .A2(n5309), .A3(n5310), .A4(n5311), .ZN(n5298)
         );
  NAND4_X1 U1646 ( .A1(n5300), .A2(n5301), .A3(n5302), .A4(n5303), .ZN(n5299)
         );
  OAI221_X1 U1647 ( .B1(n6073), .B2(n3024), .C1(n1696), .C2(n5092), .A(n5221), 
        .ZN(n3077) );
  OAI21_X1 U1648 ( .B1(n5222), .B2(n5223), .A(n6276), .ZN(n5221) );
  NAND4_X1 U1649 ( .A1(n5232), .A2(n5233), .A3(n5234), .A4(n5235), .ZN(n5222)
         );
  NAND4_X1 U1650 ( .A1(n5224), .A2(n5225), .A3(n5226), .A4(n5227), .ZN(n5223)
         );
  OAI221_X1 U1651 ( .B1(n6073), .B2(n3023), .C1(n1694), .C2(n6074), .A(n5202), 
        .ZN(n3078) );
  OAI21_X1 U1652 ( .B1(n5203), .B2(n5204), .A(n6275), .ZN(n5202) );
  NAND4_X1 U1653 ( .A1(n5213), .A2(n5214), .A3(n5215), .A4(n5216), .ZN(n5203)
         );
  NAND4_X1 U1654 ( .A1(n5205), .A2(n5206), .A3(n5207), .A4(n5208), .ZN(n5204)
         );
  OAI221_X1 U1655 ( .B1(n6073), .B2(n3022), .C1(n1692), .C2(n6075), .A(n5183), 
        .ZN(n3079) );
  OAI21_X1 U1656 ( .B1(n5184), .B2(n5185), .A(n6276), .ZN(n5183) );
  NAND4_X1 U1657 ( .A1(n5194), .A2(n5195), .A3(n5196), .A4(n5197), .ZN(n5184)
         );
  NAND4_X1 U1658 ( .A1(n5186), .A2(n5187), .A3(n5188), .A4(n5189), .ZN(n5185)
         );
  OAI221_X1 U1659 ( .B1(n5091), .B2(n3021), .C1(n1690), .C2(n5092), .A(n5164), 
        .ZN(n3080) );
  OAI21_X1 U1660 ( .B1(n5165), .B2(n5166), .A(n6274), .ZN(n5164) );
  NAND4_X1 U1661 ( .A1(n5175), .A2(n5176), .A3(n5177), .A4(n5178), .ZN(n5165)
         );
  NAND4_X1 U1662 ( .A1(n5167), .A2(n5168), .A3(n5169), .A4(n5170), .ZN(n5166)
         );
  OAI221_X1 U1663 ( .B1(n5091), .B2(n3020), .C1(n1688), .C2(n6074), .A(n5145), 
        .ZN(n3081) );
  OAI21_X1 U1664 ( .B1(n5146), .B2(n5147), .A(n6274), .ZN(n5145) );
  NAND4_X1 U1665 ( .A1(n5156), .A2(n5157), .A3(n5158), .A4(n5159), .ZN(n5146)
         );
  NAND4_X1 U1666 ( .A1(n5148), .A2(n5149), .A3(n5150), .A4(n5151), .ZN(n5147)
         );
  OAI221_X1 U1667 ( .B1(n5091), .B2(n3019), .C1(n1685), .C2(n6075), .A(n5093), 
        .ZN(n3082) );
  OAI21_X1 U1668 ( .B1(n5094), .B2(n5095), .A(n6275), .ZN(n5093) );
  NAND4_X1 U1669 ( .A1(n5121), .A2(n5122), .A3(n5123), .A4(n5124), .ZN(n5094)
         );
  NAND4_X1 U1670 ( .A1(n5097), .A2(n5098), .A3(n5099), .A4(n5100), .ZN(n5095)
         );
  OAI221_X1 U1671 ( .B1(n6278), .B2(n3018), .C1(n1748), .C2(n6279), .A(n5047), 
        .ZN(n3083) );
  OAI21_X1 U1672 ( .B1(n5048), .B2(n5049), .A(n6489), .ZN(n5047) );
  NAND4_X1 U1673 ( .A1(n5071), .A2(n5072), .A3(n5073), .A4(n5074), .ZN(n5048)
         );
  NAND4_X1 U1674 ( .A1(n5051), .A2(n5052), .A3(n5053), .A4(n5054), .ZN(n5049)
         );
  OAI221_X1 U1675 ( .B1(n4392), .B2(n3016), .C1(n1746), .C2(n6280), .A(n5027), 
        .ZN(n3085) );
  OAI21_X1 U1676 ( .B1(n5028), .B2(n5029), .A(n6490), .ZN(n5027) );
  NAND4_X1 U1677 ( .A1(n5038), .A2(n5039), .A3(n5040), .A4(n5041), .ZN(n5028)
         );
  NAND4_X1 U1678 ( .A1(n5030), .A2(n5031), .A3(n5032), .A4(n5033), .ZN(n5029)
         );
  OAI221_X1 U1679 ( .B1(n6278), .B2(n3012), .C1(n1742), .C2(n6279), .A(n4987), 
        .ZN(n3089) );
  OAI21_X1 U1680 ( .B1(n4988), .B2(n4989), .A(n6488), .ZN(n4987) );
  NAND4_X1 U1681 ( .A1(n4998), .A2(n4999), .A3(n5000), .A4(n5001), .ZN(n4988)
         );
  NAND4_X1 U1682 ( .A1(n4990), .A2(n4991), .A3(n4992), .A4(n4993), .ZN(n4989)
         );
  OAI221_X1 U1683 ( .B1(n4392), .B2(n3010), .C1(n1740), .C2(n6280), .A(n4967), 
        .ZN(n3091) );
  OAI21_X1 U1684 ( .B1(n4968), .B2(n4969), .A(n6489), .ZN(n4967) );
  NAND4_X1 U1685 ( .A1(n4978), .A2(n4979), .A3(n4980), .A4(n4981), .ZN(n4968)
         );
  NAND4_X1 U1686 ( .A1(n4970), .A2(n4971), .A3(n4972), .A4(n4973), .ZN(n4969)
         );
  OAI221_X1 U1687 ( .B1(n6278), .B2(n3006), .C1(n1736), .C2(n6279), .A(n4927), 
        .ZN(n3095) );
  OAI21_X1 U1688 ( .B1(n4928), .B2(n4929), .A(n6490), .ZN(n4927) );
  NAND4_X1 U1689 ( .A1(n4938), .A2(n4939), .A3(n4940), .A4(n4941), .ZN(n4928)
         );
  NAND4_X1 U1690 ( .A1(n4930), .A2(n4931), .A3(n4932), .A4(n4933), .ZN(n4929)
         );
  OAI221_X1 U1691 ( .B1(n4392), .B2(n3004), .C1(n1734), .C2(n6280), .A(n4907), 
        .ZN(n3097) );
  OAI21_X1 U1692 ( .B1(n4908), .B2(n4909), .A(n6488), .ZN(n4907) );
  NAND4_X1 U1693 ( .A1(n4918), .A2(n4919), .A3(n4920), .A4(n4921), .ZN(n4908)
         );
  NAND4_X1 U1694 ( .A1(n4910), .A2(n4911), .A3(n4912), .A4(n4913), .ZN(n4909)
         );
  OAI221_X1 U1695 ( .B1(n6278), .B2(n3000), .C1(n1730), .C2(n6279), .A(n4867), 
        .ZN(n3101) );
  OAI21_X1 U1696 ( .B1(n4868), .B2(n4869), .A(n6489), .ZN(n4867) );
  NAND4_X1 U1697 ( .A1(n4878), .A2(n4879), .A3(n4880), .A4(n4881), .ZN(n4868)
         );
  NAND4_X1 U1698 ( .A1(n4870), .A2(n4871), .A3(n4872), .A4(n4873), .ZN(n4869)
         );
  OAI221_X1 U1699 ( .B1(n4392), .B2(n2998), .C1(n1728), .C2(n6280), .A(n4847), 
        .ZN(n3103) );
  OAI21_X1 U1700 ( .B1(n4848), .B2(n4849), .A(n6490), .ZN(n4847) );
  NAND4_X1 U1701 ( .A1(n4858), .A2(n4859), .A3(n4860), .A4(n4861), .ZN(n4848)
         );
  NAND4_X1 U1702 ( .A1(n4850), .A2(n4851), .A3(n4852), .A4(n4853), .ZN(n4849)
         );
  OAI221_X1 U1703 ( .B1(n6278), .B2(n2994), .C1(n1724), .C2(n6279), .A(n4807), 
        .ZN(n3107) );
  OAI21_X1 U1704 ( .B1(n4808), .B2(n4809), .A(n6488), .ZN(n4807) );
  NAND4_X1 U1705 ( .A1(n4818), .A2(n4819), .A3(n4820), .A4(n4821), .ZN(n4808)
         );
  NAND4_X1 U1706 ( .A1(n4810), .A2(n4811), .A3(n4812), .A4(n4813), .ZN(n4809)
         );
  OAI221_X1 U1707 ( .B1(n4392), .B2(n2992), .C1(n1722), .C2(n6280), .A(n4787), 
        .ZN(n3109) );
  OAI21_X1 U1708 ( .B1(n4788), .B2(n4789), .A(n6489), .ZN(n4787) );
  NAND4_X1 U1709 ( .A1(n4798), .A2(n4799), .A3(n4800), .A4(n4801), .ZN(n4788)
         );
  NAND4_X1 U1710 ( .A1(n4790), .A2(n4791), .A3(n4792), .A4(n4793), .ZN(n4789)
         );
  OAI221_X1 U1711 ( .B1(n6278), .B2(n2988), .C1(n1718), .C2(n6279), .A(n4747), 
        .ZN(n3113) );
  OAI21_X1 U1712 ( .B1(n4748), .B2(n4749), .A(n6490), .ZN(n4747) );
  NAND4_X1 U1713 ( .A1(n4758), .A2(n4759), .A3(n4760), .A4(n4761), .ZN(n4748)
         );
  NAND4_X1 U1714 ( .A1(n4750), .A2(n4751), .A3(n4752), .A4(n4753), .ZN(n4749)
         );
  OAI221_X1 U1715 ( .B1(n4392), .B2(n2986), .C1(n1716), .C2(n6280), .A(n4727), 
        .ZN(n3115) );
  OAI21_X1 U1716 ( .B1(n4728), .B2(n4729), .A(n6488), .ZN(n4727) );
  NAND4_X1 U1717 ( .A1(n4738), .A2(n4739), .A3(n4740), .A4(n4741), .ZN(n4728)
         );
  NAND4_X1 U1718 ( .A1(n4730), .A2(n4731), .A3(n4732), .A4(n4733), .ZN(n4729)
         );
  OAI221_X1 U1719 ( .B1(n6278), .B2(n2982), .C1(n1712), .C2(n6279), .A(n4687), 
        .ZN(n3119) );
  OAI21_X1 U1720 ( .B1(n4688), .B2(n4689), .A(n6489), .ZN(n4687) );
  NAND4_X1 U1721 ( .A1(n4698), .A2(n4699), .A3(n4700), .A4(n4701), .ZN(n4688)
         );
  NAND4_X1 U1722 ( .A1(n4690), .A2(n4691), .A3(n4692), .A4(n4693), .ZN(n4689)
         );
  OAI221_X1 U1723 ( .B1(n4392), .B2(n2980), .C1(n1710), .C2(n6280), .A(n4667), 
        .ZN(n3121) );
  OAI21_X1 U1724 ( .B1(n4668), .B2(n4669), .A(n6490), .ZN(n4667) );
  NAND4_X1 U1725 ( .A1(n4678), .A2(n4679), .A3(n4680), .A4(n4681), .ZN(n4668)
         );
  NAND4_X1 U1726 ( .A1(n4670), .A2(n4671), .A3(n4672), .A4(n4673), .ZN(n4669)
         );
  OAI221_X1 U1727 ( .B1(n6278), .B2(n2976), .C1(n1706), .C2(n6279), .A(n4627), 
        .ZN(n3125) );
  OAI21_X1 U1728 ( .B1(n4628), .B2(n4629), .A(n6488), .ZN(n4627) );
  NAND4_X1 U1729 ( .A1(n4638), .A2(n4639), .A3(n4640), .A4(n4641), .ZN(n4628)
         );
  NAND4_X1 U1730 ( .A1(n4630), .A2(n4631), .A3(n4632), .A4(n4633), .ZN(n4629)
         );
  OAI221_X1 U1731 ( .B1(n4392), .B2(n2974), .C1(n1704), .C2(n6280), .A(n4607), 
        .ZN(n3127) );
  OAI21_X1 U1732 ( .B1(n4608), .B2(n4609), .A(n6489), .ZN(n4607) );
  NAND4_X1 U1733 ( .A1(n4618), .A2(n4619), .A3(n4620), .A4(n4621), .ZN(n4608)
         );
  NAND4_X1 U1734 ( .A1(n4610), .A2(n4611), .A3(n4612), .A4(n4613), .ZN(n4609)
         );
  OAI221_X1 U1735 ( .B1(n6278), .B2(n2966), .C1(n1696), .C2(n4393), .A(n4527), 
        .ZN(n3135) );
  OAI21_X1 U1736 ( .B1(n4528), .B2(n4529), .A(n6490), .ZN(n4527) );
  NAND4_X1 U1737 ( .A1(n4538), .A2(n4539), .A3(n4540), .A4(n4541), .ZN(n4528)
         );
  NAND4_X1 U1738 ( .A1(n4530), .A2(n4531), .A3(n4532), .A4(n4533), .ZN(n4529)
         );
  OAI221_X1 U1739 ( .B1(n6278), .B2(n2964), .C1(n1694), .C2(n6279), .A(n4507), 
        .ZN(n3137) );
  OAI21_X1 U1740 ( .B1(n4508), .B2(n4509), .A(n6489), .ZN(n4507) );
  NAND4_X1 U1741 ( .A1(n4518), .A2(n4519), .A3(n4520), .A4(n4521), .ZN(n4508)
         );
  NAND4_X1 U1742 ( .A1(n4510), .A2(n4511), .A3(n4512), .A4(n4513), .ZN(n4509)
         );
  OAI221_X1 U1743 ( .B1(n6278), .B2(n2962), .C1(n1692), .C2(n6280), .A(n4487), 
        .ZN(n3139) );
  OAI21_X1 U1744 ( .B1(n4488), .B2(n4489), .A(n6490), .ZN(n4487) );
  NAND4_X1 U1745 ( .A1(n4498), .A2(n4499), .A3(n4500), .A4(n4501), .ZN(n4488)
         );
  NAND4_X1 U1746 ( .A1(n4490), .A2(n4491), .A3(n4492), .A4(n4493), .ZN(n4489)
         );
  OAI221_X1 U1747 ( .B1(n4392), .B2(n2960), .C1(n1690), .C2(n4393), .A(n4467), 
        .ZN(n3141) );
  OAI21_X1 U1748 ( .B1(n4468), .B2(n4469), .A(n6488), .ZN(n4467) );
  NAND4_X1 U1749 ( .A1(n4478), .A2(n4479), .A3(n4480), .A4(n4481), .ZN(n4468)
         );
  NAND4_X1 U1750 ( .A1(n4470), .A2(n4471), .A3(n4472), .A4(n4473), .ZN(n4469)
         );
  OAI221_X1 U1751 ( .B1(n4392), .B2(n2958), .C1(n1688), .C2(n6279), .A(n4447), 
        .ZN(n3143) );
  OAI21_X1 U1752 ( .B1(n4448), .B2(n4449), .A(n6488), .ZN(n4447) );
  NAND4_X1 U1753 ( .A1(n4458), .A2(n4459), .A3(n4460), .A4(n4461), .ZN(n4448)
         );
  NAND4_X1 U1754 ( .A1(n4450), .A2(n4451), .A3(n4452), .A4(n4453), .ZN(n4449)
         );
  OAI221_X1 U1755 ( .B1(n4392), .B2(n2956), .C1(n1685), .C2(n6280), .A(n4394), 
        .ZN(n3145) );
  OAI21_X1 U1756 ( .B1(n4395), .B2(n4396), .A(n6489), .ZN(n4394) );
  NAND4_X1 U1757 ( .A1(n4422), .A2(n4423), .A3(n4424), .A4(n4425), .ZN(n4395)
         );
  NAND4_X1 U1758 ( .A1(n4398), .A2(n4399), .A3(n4400), .A4(n4401), .ZN(n4396)
         );
  OAI221_X1 U1759 ( .B1(n6072), .B2(n3048), .C1(n1744), .C2(n5092), .A(n5677), 
        .ZN(n3053) );
  OAI21_X1 U1760 ( .B1(n5678), .B2(n5679), .A(n6274), .ZN(n5677) );
  NAND4_X1 U1761 ( .A1(n5688), .A2(n5689), .A3(n5690), .A4(n5691), .ZN(n5678)
         );
  NAND4_X1 U1762 ( .A1(n5680), .A2(n5681), .A3(n5682), .A4(n5683), .ZN(n5679)
         );
  OAI221_X1 U1763 ( .B1(n6072), .B2(n3045), .C1(n1738), .C2(n5092), .A(n5620), 
        .ZN(n3056) );
  OAI21_X1 U1764 ( .B1(n5621), .B2(n5622), .A(n6275), .ZN(n5620) );
  NAND4_X1 U1765 ( .A1(n5631), .A2(n5632), .A3(n5633), .A4(n5634), .ZN(n5621)
         );
  NAND4_X1 U1766 ( .A1(n5623), .A2(n5624), .A3(n5625), .A4(n5626), .ZN(n5622)
         );
  OAI221_X1 U1767 ( .B1(n6072), .B2(n3042), .C1(n1732), .C2(n5092), .A(n5563), 
        .ZN(n3059) );
  OAI21_X1 U1768 ( .B1(n5564), .B2(n5565), .A(n6276), .ZN(n5563) );
  NAND4_X1 U1769 ( .A1(n5574), .A2(n5575), .A3(n5576), .A4(n5577), .ZN(n5564)
         );
  NAND4_X1 U1770 ( .A1(n5566), .A2(n5567), .A3(n5568), .A4(n5569), .ZN(n5565)
         );
  OAI221_X1 U1771 ( .B1(n6072), .B2(n3039), .C1(n1726), .C2(n5092), .A(n5506), 
        .ZN(n3062) );
  OAI21_X1 U1772 ( .B1(n5507), .B2(n5508), .A(n6274), .ZN(n5506) );
  NAND4_X1 U1773 ( .A1(n5517), .A2(n5518), .A3(n5519), .A4(n5520), .ZN(n5507)
         );
  NAND4_X1 U1774 ( .A1(n5509), .A2(n5510), .A3(n5511), .A4(n5512), .ZN(n5508)
         );
  OAI221_X1 U1775 ( .B1(n6072), .B2(n3036), .C1(n1720), .C2(n5092), .A(n5449), 
        .ZN(n3065) );
  OAI21_X1 U1776 ( .B1(n5450), .B2(n5451), .A(n6275), .ZN(n5449) );
  NAND4_X1 U1777 ( .A1(n5460), .A2(n5461), .A3(n5462), .A4(n5463), .ZN(n5450)
         );
  NAND4_X1 U1778 ( .A1(n5452), .A2(n5453), .A3(n5454), .A4(n5455), .ZN(n5451)
         );
  OAI221_X1 U1779 ( .B1(n6072), .B2(n3033), .C1(n1714), .C2(n5092), .A(n5392), 
        .ZN(n3068) );
  OAI21_X1 U1780 ( .B1(n5393), .B2(n5394), .A(n6276), .ZN(n5392) );
  NAND4_X1 U1781 ( .A1(n5403), .A2(n5404), .A3(n5405), .A4(n5406), .ZN(n5393)
         );
  NAND4_X1 U1782 ( .A1(n5395), .A2(n5396), .A3(n5397), .A4(n5398), .ZN(n5394)
         );
  OAI221_X1 U1783 ( .B1(n6072), .B2(n3030), .C1(n1708), .C2(n5092), .A(n5335), 
        .ZN(n3071) );
  OAI21_X1 U1784 ( .B1(n5336), .B2(n5337), .A(n6274), .ZN(n5335) );
  NAND4_X1 U1785 ( .A1(n5346), .A2(n5347), .A3(n5348), .A4(n5349), .ZN(n5336)
         );
  NAND4_X1 U1786 ( .A1(n5338), .A2(n5339), .A3(n5340), .A4(n5341), .ZN(n5337)
         );
  OAI221_X1 U1787 ( .B1(n6072), .B2(n3027), .C1(n1702), .C2(n5092), .A(n5278), 
        .ZN(n3074) );
  OAI21_X1 U1788 ( .B1(n5279), .B2(n5280), .A(n6275), .ZN(n5278) );
  NAND4_X1 U1789 ( .A1(n5289), .A2(n5290), .A3(n5291), .A4(n5292), .ZN(n5279)
         );
  NAND4_X1 U1790 ( .A1(n5281), .A2(n5282), .A3(n5283), .A4(n5284), .ZN(n5280)
         );
  OAI221_X1 U1791 ( .B1(n6072), .B2(n3026), .C1(n1700), .C2(n6074), .A(n5259), 
        .ZN(n3075) );
  OAI21_X1 U1792 ( .B1(n5260), .B2(n5261), .A(n6276), .ZN(n5259) );
  NAND4_X1 U1793 ( .A1(n5270), .A2(n5271), .A3(n5272), .A4(n5273), .ZN(n5260)
         );
  NAND4_X1 U1794 ( .A1(n5262), .A2(n5263), .A3(n5264), .A4(n5265), .ZN(n5261)
         );
  OAI221_X1 U1795 ( .B1(n6072), .B2(n3025), .C1(n1698), .C2(n6075), .A(n5240), 
        .ZN(n3076) );
  OAI21_X1 U1796 ( .B1(n5241), .B2(n5242), .A(n6274), .ZN(n5240) );
  NAND4_X1 U1797 ( .A1(n5251), .A2(n5252), .A3(n5253), .A4(n5254), .ZN(n5241)
         );
  NAND4_X1 U1798 ( .A1(n5243), .A2(n5244), .A3(n5245), .A4(n5246), .ZN(n5242)
         );
  OAI221_X1 U1799 ( .B1(n6277), .B2(n3014), .C1(n1744), .C2(n4393), .A(n5007), 
        .ZN(n3087) );
  OAI21_X1 U1800 ( .B1(n5008), .B2(n5009), .A(n6488), .ZN(n5007) );
  NAND4_X1 U1801 ( .A1(n5018), .A2(n5019), .A3(n5020), .A4(n5021), .ZN(n5008)
         );
  NAND4_X1 U1802 ( .A1(n5010), .A2(n5011), .A3(n5012), .A4(n5013), .ZN(n5009)
         );
  OAI221_X1 U1803 ( .B1(n6277), .B2(n3008), .C1(n1738), .C2(n4393), .A(n4947), 
        .ZN(n3093) );
  OAI21_X1 U1804 ( .B1(n4948), .B2(n4949), .A(n6489), .ZN(n4947) );
  NAND4_X1 U1805 ( .A1(n4958), .A2(n4959), .A3(n4960), .A4(n4961), .ZN(n4948)
         );
  NAND4_X1 U1806 ( .A1(n4950), .A2(n4951), .A3(n4952), .A4(n4953), .ZN(n4949)
         );
  OAI221_X1 U1807 ( .B1(n6277), .B2(n3002), .C1(n1732), .C2(n4393), .A(n4887), 
        .ZN(n3099) );
  OAI21_X1 U1808 ( .B1(n4888), .B2(n4889), .A(n6490), .ZN(n4887) );
  NAND4_X1 U1809 ( .A1(n4898), .A2(n4899), .A3(n4900), .A4(n4901), .ZN(n4888)
         );
  NAND4_X1 U1810 ( .A1(n4890), .A2(n4891), .A3(n4892), .A4(n4893), .ZN(n4889)
         );
  OAI221_X1 U1811 ( .B1(n6277), .B2(n2996), .C1(n1726), .C2(n4393), .A(n4827), 
        .ZN(n3105) );
  OAI21_X1 U1812 ( .B1(n4828), .B2(n4829), .A(n6488), .ZN(n4827) );
  NAND4_X1 U1813 ( .A1(n4838), .A2(n4839), .A3(n4840), .A4(n4841), .ZN(n4828)
         );
  NAND4_X1 U1814 ( .A1(n4830), .A2(n4831), .A3(n4832), .A4(n4833), .ZN(n4829)
         );
  OAI221_X1 U1815 ( .B1(n6277), .B2(n2990), .C1(n1720), .C2(n4393), .A(n4767), 
        .ZN(n3111) );
  OAI21_X1 U1816 ( .B1(n4768), .B2(n4769), .A(n6489), .ZN(n4767) );
  NAND4_X1 U1817 ( .A1(n4778), .A2(n4779), .A3(n4780), .A4(n4781), .ZN(n4768)
         );
  NAND4_X1 U1818 ( .A1(n4770), .A2(n4771), .A3(n4772), .A4(n4773), .ZN(n4769)
         );
  OAI221_X1 U1819 ( .B1(n6277), .B2(n2984), .C1(n1714), .C2(n4393), .A(n4707), 
        .ZN(n3117) );
  OAI21_X1 U1820 ( .B1(n4708), .B2(n4709), .A(n6490), .ZN(n4707) );
  NAND4_X1 U1821 ( .A1(n4718), .A2(n4719), .A3(n4720), .A4(n4721), .ZN(n4708)
         );
  NAND4_X1 U1822 ( .A1(n4710), .A2(n4711), .A3(n4712), .A4(n4713), .ZN(n4709)
         );
  OAI221_X1 U1823 ( .B1(n6277), .B2(n2978), .C1(n1708), .C2(n4393), .A(n4647), 
        .ZN(n3123) );
  OAI21_X1 U1824 ( .B1(n4648), .B2(n4649), .A(n6488), .ZN(n4647) );
  NAND4_X1 U1825 ( .A1(n4658), .A2(n4659), .A3(n4660), .A4(n4661), .ZN(n4648)
         );
  NAND4_X1 U1826 ( .A1(n4650), .A2(n4651), .A3(n4652), .A4(n4653), .ZN(n4649)
         );
  OAI221_X1 U1827 ( .B1(n6277), .B2(n2972), .C1(n1702), .C2(n4393), .A(n4587), 
        .ZN(n3129) );
  OAI21_X1 U1828 ( .B1(n4588), .B2(n4589), .A(n6489), .ZN(n4587) );
  NAND4_X1 U1829 ( .A1(n4598), .A2(n4599), .A3(n4600), .A4(n4601), .ZN(n4588)
         );
  NAND4_X1 U1830 ( .A1(n4590), .A2(n4591), .A3(n4592), .A4(n4593), .ZN(n4589)
         );
  OAI221_X1 U1831 ( .B1(n6277), .B2(n2970), .C1(n1700), .C2(n6279), .A(n4567), 
        .ZN(n3131) );
  OAI21_X1 U1832 ( .B1(n4568), .B2(n4569), .A(n6490), .ZN(n4567) );
  NAND4_X1 U1833 ( .A1(n4578), .A2(n4579), .A3(n4580), .A4(n4581), .ZN(n4568)
         );
  NAND4_X1 U1834 ( .A1(n4570), .A2(n4571), .A3(n4572), .A4(n4573), .ZN(n4569)
         );
  OAI221_X1 U1835 ( .B1(n6277), .B2(n2968), .C1(n1698), .C2(n6280), .A(n4547), 
        .ZN(n3133) );
  OAI21_X1 U1836 ( .B1(n4548), .B2(n4549), .A(n6488), .ZN(n4547) );
  NAND4_X1 U1837 ( .A1(n4558), .A2(n4559), .A3(n4560), .A4(n4561), .ZN(n4548)
         );
  NAND4_X1 U1838 ( .A1(n4550), .A2(n4551), .A3(n4552), .A4(n4553), .ZN(n4549)
         );
  AOI221_X1 U1839 ( .B1(n6235), .B2(\registers[13][0] ), .C1(n6243), .C2(
        \registers[12][0] ), .A(n5728), .ZN(n5721) );
  OAI22_X1 U1840 ( .A1(n2792), .A2(n6247), .B1(n5784), .B2(n6260), .ZN(n5728)
         );
  AOI221_X1 U1841 ( .B1(n6182), .B2(\registers[31][0] ), .C1(n6184), .C2(
        \registers[30][0] ), .A(n5734), .ZN(n5719) );
  OAI22_X1 U1842 ( .A1(n2852), .A2(n6187), .B1(n5842), .B2(n6195), .ZN(n5734)
         );
  AOI221_X1 U1843 ( .B1(n6203), .B2(\registers[21][0] ), .C1(n6214), .C2(
        \registers[20][0] ), .A(n5731), .ZN(n5720) );
  OAI22_X1 U1844 ( .A1(n2793), .A2(n6219), .B1(n5785), .B2(n6227), .ZN(n5731)
         );
  AOI221_X1 U1845 ( .B1(n6109), .B2(\registers[29][0] ), .C1(n6117), .C2(
        \registers[28][0] ), .A(n5747), .ZN(n5740) );
  OAI22_X1 U1846 ( .A1(n4220), .A2(n6125), .B1(n5918), .B2(n6129), .ZN(n5747)
         );
  AOI221_X1 U1847 ( .B1(n6077), .B2(\registers[23][0] ), .C1(n6088), .C2(
        \registers[22][0] ), .A(n5750), .ZN(n5739) );
  OAI22_X1 U1848 ( .A1(n2853), .A2(n6096), .B1(n5843), .B2(n6107), .ZN(n5750)
         );
  AOI221_X1 U1849 ( .B1(n6236), .B2(\registers[13][1] ), .C1(n6244), .C2(
        \registers[12][1] ), .A(n5704), .ZN(n5701) );
  OAI22_X1 U1850 ( .A1(n2794), .A2(n6251), .B1(n5786), .B2(n6259), .ZN(n5704)
         );
  AOI221_X1 U1851 ( .B1(n6183), .B2(\registers[31][1] ), .C1(n6185), .C2(
        \registers[30][1] ), .A(n5706), .ZN(n5699) );
  OAI22_X1 U1852 ( .A1(n2854), .A2(n6190), .B1(n5844), .B2(n6197), .ZN(n5706)
         );
  AOI221_X1 U1853 ( .B1(n6204), .B2(\registers[21][1] ), .C1(n6211), .C2(
        \registers[20][1] ), .A(n5705), .ZN(n5700) );
  OAI22_X1 U1854 ( .A1(n2795), .A2(n6222), .B1(n5787), .B2(n6230), .ZN(n5705)
         );
  AOI221_X1 U1855 ( .B1(n6115), .B2(\registers[29][1] ), .C1(n6118), .C2(
        \registers[28][1] ), .A(n5713), .ZN(n5708) );
  OAI22_X1 U1856 ( .A1(n4221), .A2(n6121), .B1(n5919), .B2(n6131), .ZN(n5713)
         );
  AOI221_X1 U1857 ( .B1(n6078), .B2(\registers[23][1] ), .C1(n6088), .C2(
        \registers[22][1] ), .A(n5714), .ZN(n5707) );
  OAI22_X1 U1858 ( .A1(n2855), .A2(n6093), .B1(n5845), .B2(n6101), .ZN(n5714)
         );
  AOI221_X1 U1859 ( .B1(n6236), .B2(\registers[13][2] ), .C1(n6242), .C2(
        \registers[12][2] ), .A(n5685), .ZN(n5682) );
  OAI22_X1 U1860 ( .A1(n2796), .A2(n6251), .B1(n5788), .B2(n6259), .ZN(n5685)
         );
  AOI221_X1 U1861 ( .B1(n5116), .B2(\registers[31][2] ), .C1(n5117), .C2(
        \registers[30][2] ), .A(n5687), .ZN(n5680) );
  OAI22_X1 U1862 ( .A1(n2856), .A2(n6193), .B1(n5846), .B2(n6199), .ZN(n5687)
         );
  AOI221_X1 U1863 ( .B1(n6204), .B2(\registers[21][2] ), .C1(n6211), .C2(
        \registers[20][2] ), .A(n5686), .ZN(n5681) );
  OAI22_X1 U1864 ( .A1(n2797), .A2(n6219), .B1(n5789), .B2(n6232), .ZN(n5686)
         );
  AOI221_X1 U1865 ( .B1(n6109), .B2(\registers[29][2] ), .C1(n6116), .C2(
        \registers[28][2] ), .A(n5694), .ZN(n5689) );
  OAI22_X1 U1866 ( .A1(n4222), .A2(n6126), .B1(n5920), .B2(n6134), .ZN(n5694)
         );
  AOI221_X1 U1867 ( .B1(n6077), .B2(\registers[23][2] ), .C1(n6085), .C2(
        \registers[22][2] ), .A(n5695), .ZN(n5688) );
  OAI22_X1 U1868 ( .A1(n2857), .A2(n6098), .B1(n5847), .B2(n6106), .ZN(n5695)
         );
  AOI221_X1 U1869 ( .B1(n6237), .B2(\registers[13][3] ), .C1(n6242), .C2(
        \registers[12][3] ), .A(n5666), .ZN(n5663) );
  OAI22_X1 U1870 ( .A1(n2798), .A2(n6250), .B1(n5790), .B2(n6258), .ZN(n5666)
         );
  AOI221_X1 U1871 ( .B1(n6182), .B2(\registers[31][3] ), .C1(n6184), .C2(
        \registers[30][3] ), .A(n5668), .ZN(n5661) );
  OAI22_X1 U1872 ( .A1(n2860), .A2(n6187), .B1(n5848), .B2(n6201), .ZN(n5668)
         );
  AOI221_X1 U1873 ( .B1(n6205), .B2(\registers[21][3] ), .C1(n6212), .C2(
        \registers[20][3] ), .A(n5667), .ZN(n5662) );
  OAI22_X1 U1874 ( .A1(n2799), .A2(n6220), .B1(n5791), .B2(n6227), .ZN(n5667)
         );
  AOI221_X1 U1875 ( .B1(n6111), .B2(\registers[29][3] ), .C1(n6116), .C2(
        \registers[28][3] ), .A(n5675), .ZN(n5670) );
  OAI22_X1 U1876 ( .A1(n4223), .A2(n6124), .B1(n5921), .B2(n6132), .ZN(n5675)
         );
  AOI221_X1 U1877 ( .B1(n6079), .B2(\registers[23][3] ), .C1(n6086), .C2(
        \registers[22][3] ), .A(n5676), .ZN(n5669) );
  OAI22_X1 U1878 ( .A1(n2895), .A2(n6093), .B1(n5849), .B2(n6105), .ZN(n5676)
         );
  AOI221_X1 U1879 ( .B1(n6238), .B2(\registers[13][4] ), .C1(n6243), .C2(
        \registers[12][4] ), .A(n5647), .ZN(n5644) );
  OAI22_X1 U1880 ( .A1(n2800), .A2(n6246), .B1(n5792), .B2(n6254), .ZN(n5647)
         );
  AOI221_X1 U1881 ( .B1(n6183), .B2(\registers[31][4] ), .C1(n6185), .C2(
        \registers[30][4] ), .A(n5649), .ZN(n5642) );
  OAI22_X1 U1882 ( .A1(n2929), .A2(n6188), .B1(n5850), .B2(n6195), .ZN(n5649)
         );
  AOI221_X1 U1883 ( .B1(n6206), .B2(\registers[21][4] ), .C1(n6217), .C2(
        \registers[20][4] ), .A(n5648), .ZN(n5643) );
  OAI22_X1 U1884 ( .A1(n2801), .A2(n6220), .B1(n5793), .B2(n6228), .ZN(n5648)
         );
  AOI221_X1 U1885 ( .B1(n6112), .B2(\registers[29][4] ), .C1(n6117), .C2(
        \registers[28][4] ), .A(n5656), .ZN(n5651) );
  OAI22_X1 U1886 ( .A1(n4224), .A2(n6120), .B1(n5922), .B2(n6128), .ZN(n5656)
         );
  AOI221_X1 U1887 ( .B1(n6080), .B2(\registers[23][4] ), .C1(n6086), .C2(
        \registers[22][4] ), .A(n5657), .ZN(n5650) );
  OAI22_X1 U1888 ( .A1(n2971), .A2(n6093), .B1(n5851), .B2(n6101), .ZN(n5657)
         );
  AOI221_X1 U1889 ( .B1(n6237), .B2(\registers[13][5] ), .C1(n6243), .C2(
        \registers[12][5] ), .A(n5628), .ZN(n5625) );
  OAI22_X1 U1890 ( .A1(n2802), .A2(n6247), .B1(n5794), .B2(n6255), .ZN(n5628)
         );
  AOI221_X1 U1891 ( .B1(n5116), .B2(\registers[31][5] ), .C1(n5117), .C2(
        \registers[30][5] ), .A(n5630), .ZN(n5623) );
  OAI22_X1 U1892 ( .A1(n4150), .A2(n6189), .B1(n5852), .B2(n6196), .ZN(n5630)
         );
  AOI221_X1 U1893 ( .B1(n6203), .B2(\registers[21][5] ), .C1(n6212), .C2(
        \registers[20][5] ), .A(n5629), .ZN(n5624) );
  OAI22_X1 U1894 ( .A1(n2803), .A2(n6221), .B1(n5795), .B2(n6229), .ZN(n5629)
         );
  AOI221_X1 U1895 ( .B1(n6109), .B2(\registers[29][5] ), .C1(n6117), .C2(
        \registers[28][5] ), .A(n5637), .ZN(n5632) );
  OAI22_X1 U1896 ( .A1(n4225), .A2(n6121), .B1(n5923), .B2(n6129), .ZN(n5637)
         );
  AOI221_X1 U1897 ( .B1(n6079), .B2(\registers[23][5] ), .C1(n6090), .C2(
        \registers[22][5] ), .A(n5638), .ZN(n5631) );
  OAI22_X1 U1898 ( .A1(n4151), .A2(n6094), .B1(n5853), .B2(n6102), .ZN(n5638)
         );
  AOI221_X1 U1899 ( .B1(n6241), .B2(\registers[13][6] ), .C1(n6244), .C2(
        \registers[12][6] ), .A(n5609), .ZN(n5606) );
  OAI22_X1 U1900 ( .A1(n2804), .A2(n6248), .B1(n5796), .B2(n6257), .ZN(n5609)
         );
  AOI221_X1 U1901 ( .B1(n6182), .B2(\registers[31][6] ), .C1(n6184), .C2(
        \registers[30][6] ), .A(n5611), .ZN(n5604) );
  OAI22_X1 U1902 ( .A1(n4152), .A2(n6190), .B1(n5854), .B2(n6197), .ZN(n5611)
         );
  AOI221_X1 U1903 ( .B1(n6205), .B2(\registers[21][6] ), .C1(n6213), .C2(
        \registers[20][6] ), .A(n5610), .ZN(n5605) );
  OAI22_X1 U1904 ( .A1(n2805), .A2(n6222), .B1(n5797), .B2(n6230), .ZN(n5610)
         );
  AOI221_X1 U1905 ( .B1(n6110), .B2(\registers[29][6] ), .C1(n6118), .C2(
        \registers[28][6] ), .A(n5618), .ZN(n5613) );
  OAI22_X1 U1906 ( .A1(n4226), .A2(n6122), .B1(n5924), .B2(n6130), .ZN(n5618)
         );
  AOI221_X1 U1907 ( .B1(n6083), .B2(\registers[23][6] ), .C1(n6087), .C2(
        \registers[22][6] ), .A(n5619), .ZN(n5612) );
  OAI22_X1 U1908 ( .A1(n4153), .A2(n6095), .B1(n5855), .B2(n6103), .ZN(n5619)
         );
  AOI221_X1 U1909 ( .B1(n6239), .B2(\registers[13][7] ), .C1(n6242), .C2(
        \registers[12][7] ), .A(n5590), .ZN(n5587) );
  OAI22_X1 U1910 ( .A1(n2806), .A2(n6249), .B1(n5798), .B2(n6256), .ZN(n5590)
         );
  AOI221_X1 U1911 ( .B1(n6183), .B2(\registers[31][7] ), .C1(n6185), .C2(
        \registers[30][7] ), .A(n5592), .ZN(n5585) );
  OAI22_X1 U1912 ( .A1(n4154), .A2(n6191), .B1(n5856), .B2(n6198), .ZN(n5592)
         );
  AOI221_X1 U1913 ( .B1(n6208), .B2(\registers[21][7] ), .C1(n6214), .C2(
        \registers[20][7] ), .A(n5591), .ZN(n5586) );
  OAI22_X1 U1914 ( .A1(n2807), .A2(n6223), .B1(n5799), .B2(n6231), .ZN(n5591)
         );
  AOI221_X1 U1915 ( .B1(n6111), .B2(\registers[29][7] ), .C1(n6116), .C2(
        \registers[28][7] ), .A(n5599), .ZN(n5594) );
  OAI22_X1 U1916 ( .A1(n4227), .A2(n6123), .B1(n5925), .B2(n6129), .ZN(n5599)
         );
  AOI221_X1 U1917 ( .B1(n6081), .B2(\registers[23][7] ), .C1(n6087), .C2(
        \registers[22][7] ), .A(n5600), .ZN(n5593) );
  OAI22_X1 U1918 ( .A1(n4155), .A2(n6096), .B1(n5857), .B2(n6104), .ZN(n5600)
         );
  AOI221_X1 U1919 ( .B1(n6239), .B2(\registers[13][8] ), .C1(n6244), .C2(
        \registers[12][8] ), .A(n5571), .ZN(n5568) );
  OAI22_X1 U1920 ( .A1(n2808), .A2(n6248), .B1(n5800), .B2(n6257), .ZN(n5571)
         );
  AOI221_X1 U1921 ( .B1(n5116), .B2(\registers[31][8] ), .C1(n5117), .C2(
        \registers[30][8] ), .A(n5573), .ZN(n5566) );
  OAI22_X1 U1922 ( .A1(n4156), .A2(n6190), .B1(n5858), .B2(n6197), .ZN(n5573)
         );
  AOI221_X1 U1923 ( .B1(n6205), .B2(\registers[21][8] ), .C1(n6214), .C2(
        \registers[20][8] ), .A(n5572), .ZN(n5567) );
  OAI22_X1 U1924 ( .A1(n2809), .A2(n6222), .B1(n5801), .B2(n6230), .ZN(n5572)
         );
  AOI221_X1 U1925 ( .B1(n6110), .B2(\registers[29][8] ), .C1(n6118), .C2(
        \registers[28][8] ), .A(n5580), .ZN(n5575) );
  OAI22_X1 U1926 ( .A1(n4228), .A2(n6123), .B1(n5926), .B2(n6131), .ZN(n5580)
         );
  AOI221_X1 U1927 ( .B1(n6081), .B2(\registers[23][8] ), .C1(n6089), .C2(
        \registers[22][8] ), .A(n5581), .ZN(n5574) );
  OAI22_X1 U1928 ( .A1(n4157), .A2(n6094), .B1(n5859), .B2(n6102), .ZN(n5581)
         );
  AOI221_X1 U1929 ( .B1(n6239), .B2(\registers[13][9] ), .C1(n6243), .C2(
        \registers[12][9] ), .A(n5552), .ZN(n5549) );
  OAI22_X1 U1930 ( .A1(n2810), .A2(n6247), .B1(n5802), .B2(n6257), .ZN(n5552)
         );
  AOI221_X1 U1931 ( .B1(n6182), .B2(\registers[31][9] ), .C1(n6184), .C2(
        \registers[30][9] ), .A(n5554), .ZN(n5547) );
  OAI22_X1 U1932 ( .A1(n4158), .A2(n6189), .B1(n5860), .B2(n6196), .ZN(n5554)
         );
  AOI221_X1 U1933 ( .B1(n6207), .B2(\registers[21][9] ), .C1(n6215), .C2(
        \registers[20][9] ), .A(n5553), .ZN(n5548) );
  OAI22_X1 U1934 ( .A1(n2811), .A2(n6221), .B1(n5803), .B2(n6229), .ZN(n5553)
         );
  AOI221_X1 U1935 ( .B1(n6113), .B2(\registers[29][9] ), .C1(n6117), .C2(
        \registers[28][9] ), .A(n5561), .ZN(n5556) );
  OAI22_X1 U1936 ( .A1(n4229), .A2(n6122), .B1(n5927), .B2(n6129), .ZN(n5561)
         );
  AOI221_X1 U1937 ( .B1(n6081), .B2(\registers[23][9] ), .C1(n6089), .C2(
        \registers[22][9] ), .A(n5562), .ZN(n5555) );
  OAI22_X1 U1938 ( .A1(n4159), .A2(n6094), .B1(n5861), .B2(n6104), .ZN(n5562)
         );
  AOI221_X1 U1939 ( .B1(n6238), .B2(\registers[13][10] ), .C1(n6244), .C2(
        \registers[12][10] ), .A(n5533), .ZN(n5530) );
  OAI22_X1 U1940 ( .A1(n2812), .A2(n6250), .B1(n5804), .B2(n6258), .ZN(n5533)
         );
  AOI221_X1 U1941 ( .B1(n6183), .B2(\registers[31][10] ), .C1(n6185), .C2(
        \registers[30][10] ), .A(n5535), .ZN(n5528) );
  OAI22_X1 U1942 ( .A1(n4160), .A2(n6192), .B1(n5862), .B2(n6199), .ZN(n5535)
         );
  AOI221_X1 U1943 ( .B1(n6206), .B2(\registers[21][10] ), .C1(n6215), .C2(
        \registers[20][10] ), .A(n5534), .ZN(n5529) );
  OAI22_X1 U1944 ( .A1(n2813), .A2(n6224), .B1(n5805), .B2(n6227), .ZN(n5534)
         );
  AOI221_X1 U1945 ( .B1(n6112), .B2(\registers[29][10] ), .C1(n6118), .C2(
        \registers[28][10] ), .A(n5542), .ZN(n5537) );
  OAI22_X1 U1946 ( .A1(n4230), .A2(n6124), .B1(n5928), .B2(n6132), .ZN(n5542)
         );
  AOI221_X1 U1947 ( .B1(n6080), .B2(\registers[23][10] ), .C1(n6088), .C2(
        \registers[22][10] ), .A(n5543), .ZN(n5536) );
  OAI22_X1 U1948 ( .A1(n4161), .A2(n6097), .B1(n5863), .B2(n6101), .ZN(n5543)
         );
  AOI221_X1 U1949 ( .B1(n6239), .B2(\registers[13][11] ), .C1(n6242), .C2(
        \registers[12][11] ), .A(n5514), .ZN(n5511) );
  OAI22_X1 U1950 ( .A1(n2814), .A2(n6251), .B1(n5806), .B2(n6259), .ZN(n5514)
         );
  AOI221_X1 U1951 ( .B1(n5116), .B2(\registers[31][11] ), .C1(n5117), .C2(
        \registers[30][11] ), .A(n5516), .ZN(n5509) );
  OAI22_X1 U1952 ( .A1(n4162), .A2(n6193), .B1(n5864), .B2(n6200), .ZN(n5516)
         );
  AOI221_X1 U1953 ( .B1(n6207), .B2(\registers[21][11] ), .C1(n6215), .C2(
        \registers[20][11] ), .A(n5515), .ZN(n5510) );
  OAI22_X1 U1954 ( .A1(n2815), .A2(n6225), .B1(n5807), .B2(n6232), .ZN(n5515)
         );
  AOI221_X1 U1955 ( .B1(n6113), .B2(\registers[29][11] ), .C1(n6116), .C2(
        \registers[28][11] ), .A(n5523), .ZN(n5518) );
  OAI22_X1 U1956 ( .A1(n4231), .A2(n6126), .B1(n5929), .B2(n6133), .ZN(n5523)
         );
  AOI221_X1 U1957 ( .B1(n6081), .B2(\registers[23][11] ), .C1(n6089), .C2(
        \registers[22][11] ), .A(n5524), .ZN(n5517) );
  OAI22_X1 U1958 ( .A1(n4163), .A2(n6098), .B1(n5865), .B2(n6107), .ZN(n5524)
         );
  AOI221_X1 U1959 ( .B1(n6240), .B2(\registers[13][12] ), .C1(n6242), .C2(
        \registers[12][12] ), .A(n5495), .ZN(n5492) );
  OAI22_X1 U1960 ( .A1(n2816), .A2(n6246), .B1(n5808), .B2(n6254), .ZN(n5495)
         );
  AOI221_X1 U1961 ( .B1(n6182), .B2(\registers[31][12] ), .C1(n6184), .C2(
        \registers[30][12] ), .A(n5497), .ZN(n5490) );
  OAI22_X1 U1962 ( .A1(n4164), .A2(n6188), .B1(n5866), .B2(n6195), .ZN(n5497)
         );
  AOI221_X1 U1963 ( .B1(n6208), .B2(\registers[21][12] ), .C1(n6216), .C2(
        \registers[20][12] ), .A(n5496), .ZN(n5491) );
  OAI22_X1 U1964 ( .A1(n2817), .A2(n6220), .B1(n5809), .B2(n6228), .ZN(n5496)
         );
  AOI221_X1 U1965 ( .B1(n6114), .B2(\registers[29][12] ), .C1(n6116), .C2(
        \registers[28][12] ), .A(n5504), .ZN(n5499) );
  OAI22_X1 U1966 ( .A1(n4232), .A2(n6120), .B1(n5930), .B2(n6128), .ZN(n5504)
         );
  AOI221_X1 U1967 ( .B1(n6082), .B2(\registers[23][12] ), .C1(n6090), .C2(
        \registers[22][12] ), .A(n5505), .ZN(n5498) );
  OAI22_X1 U1968 ( .A1(n4165), .A2(n6093), .B1(n5867), .B2(n6101), .ZN(n5505)
         );
  AOI221_X1 U1969 ( .B1(n6240), .B2(\registers[13][13] ), .C1(n6243), .C2(
        \registers[12][13] ), .A(n5476), .ZN(n5473) );
  OAI22_X1 U1970 ( .A1(n2818), .A2(n6247), .B1(n5810), .B2(n6255), .ZN(n5476)
         );
  AOI221_X1 U1971 ( .B1(n6183), .B2(\registers[31][13] ), .C1(n6185), .C2(
        \registers[30][13] ), .A(n5478), .ZN(n5471) );
  OAI22_X1 U1972 ( .A1(n4166), .A2(n6189), .B1(n5868), .B2(n6196), .ZN(n5478)
         );
  AOI221_X1 U1973 ( .B1(n6208), .B2(\registers[21][13] ), .C1(n6216), .C2(
        \registers[20][13] ), .A(n5477), .ZN(n5472) );
  OAI22_X1 U1974 ( .A1(n2819), .A2(n6221), .B1(n5811), .B2(n6229), .ZN(n5477)
         );
  AOI221_X1 U1975 ( .B1(n6114), .B2(\registers[29][13] ), .C1(n6117), .C2(
        \registers[28][13] ), .A(n5485), .ZN(n5480) );
  OAI22_X1 U1976 ( .A1(n4233), .A2(n6121), .B1(n5931), .B2(n6129), .ZN(n5485)
         );
  AOI221_X1 U1977 ( .B1(n6082), .B2(\registers[23][13] ), .C1(n6090), .C2(
        \registers[22][13] ), .A(n5486), .ZN(n5479) );
  OAI22_X1 U1978 ( .A1(n4167), .A2(n6094), .B1(n5869), .B2(n6102), .ZN(n5486)
         );
  AOI221_X1 U1979 ( .B1(n6238), .B2(\registers[13][14] ), .C1(n6243), .C2(
        \registers[12][14] ), .A(n5457), .ZN(n5454) );
  OAI22_X1 U1980 ( .A1(n2820), .A2(n6248), .B1(n5812), .B2(n6255), .ZN(n5457)
         );
  AOI221_X1 U1981 ( .B1(n5116), .B2(\registers[31][14] ), .C1(n5117), .C2(
        \registers[30][14] ), .A(n5459), .ZN(n5452) );
  OAI22_X1 U1982 ( .A1(n4168), .A2(n6190), .B1(n5870), .B2(n6197), .ZN(n5459)
         );
  AOI221_X1 U1983 ( .B1(n6206), .B2(\registers[21][14] ), .C1(n6215), .C2(
        \registers[20][14] ), .A(n5458), .ZN(n5453) );
  OAI22_X1 U1984 ( .A1(n2821), .A2(n6222), .B1(n5813), .B2(n6230), .ZN(n5458)
         );
  AOI221_X1 U1985 ( .B1(n6112), .B2(\registers[29][14] ), .C1(n6117), .C2(
        \registers[28][14] ), .A(n5466), .ZN(n5461) );
  OAI22_X1 U1986 ( .A1(n4234), .A2(n6122), .B1(n5932), .B2(n6130), .ZN(n5466)
         );
  AOI221_X1 U1987 ( .B1(n6080), .B2(\registers[23][14] ), .C1(n6088), .C2(
        \registers[22][14] ), .A(n5467), .ZN(n5460) );
  OAI22_X1 U1988 ( .A1(n4169), .A2(n6095), .B1(n5871), .B2(n6103), .ZN(n5467)
         );
  AOI221_X1 U1989 ( .B1(n6239), .B2(\registers[13][15] ), .C1(n6244), .C2(
        \registers[12][15] ), .A(n5438), .ZN(n5435) );
  OAI22_X1 U1990 ( .A1(n2822), .A2(n6249), .B1(n5814), .B2(n6256), .ZN(n5438)
         );
  AOI221_X1 U1991 ( .B1(n6182), .B2(\registers[31][15] ), .C1(n6184), .C2(
        \registers[30][15] ), .A(n5440), .ZN(n5433) );
  OAI22_X1 U1992 ( .A1(n4170), .A2(n6191), .B1(n5872), .B2(n6198), .ZN(n5440)
         );
  AOI221_X1 U1993 ( .B1(n6207), .B2(\registers[21][15] ), .C1(n6211), .C2(
        \registers[20][15] ), .A(n5439), .ZN(n5434) );
  OAI22_X1 U1994 ( .A1(n2823), .A2(n6223), .B1(n5815), .B2(n6231), .ZN(n5439)
         );
  AOI221_X1 U1995 ( .B1(n6113), .B2(\registers[29][15] ), .C1(n6118), .C2(
        \registers[28][15] ), .A(n5447), .ZN(n5442) );
  OAI22_X1 U1996 ( .A1(n4235), .A2(n6123), .B1(n5933), .B2(n6130), .ZN(n5447)
         );
  AOI221_X1 U1997 ( .B1(n6081), .B2(\registers[23][15] ), .C1(n6089), .C2(
        \registers[22][15] ), .A(n5448), .ZN(n5441) );
  OAI22_X1 U1998 ( .A1(n4171), .A2(n6096), .B1(n5873), .B2(n6103), .ZN(n5448)
         );
  AOI221_X1 U1999 ( .B1(n6240), .B2(\registers[13][16] ), .C1(n6242), .C2(
        \registers[12][16] ), .A(n5419), .ZN(n5416) );
  OAI22_X1 U2000 ( .A1(n2826), .A2(n6249), .B1(n5816), .B2(n6256), .ZN(n5419)
         );
  AOI221_X1 U2001 ( .B1(n6183), .B2(\registers[31][16] ), .C1(n6185), .C2(
        \registers[30][16] ), .A(n5421), .ZN(n5414) );
  OAI22_X1 U2002 ( .A1(n4172), .A2(n6191), .B1(n5874), .B2(n6198), .ZN(n5421)
         );
  AOI221_X1 U2003 ( .B1(n6208), .B2(\registers[21][16] ), .C1(n6216), .C2(
        \registers[20][16] ), .A(n5420), .ZN(n5415) );
  OAI22_X1 U2004 ( .A1(n2827), .A2(n6223), .B1(n5817), .B2(n6229), .ZN(n5420)
         );
  AOI221_X1 U2005 ( .B1(n6114), .B2(\registers[29][16] ), .C1(n6116), .C2(
        \registers[28][16] ), .A(n5428), .ZN(n5423) );
  OAI22_X1 U2006 ( .A1(n4236), .A2(n6122), .B1(n5934), .B2(n6131), .ZN(n5428)
         );
  AOI221_X1 U2007 ( .B1(n6082), .B2(\registers[23][16] ), .C1(n6090), .C2(
        \registers[22][16] ), .A(n5429), .ZN(n5422) );
  OAI22_X1 U2008 ( .A1(n4173), .A2(n6095), .B1(n5875), .B2(n6104), .ZN(n5429)
         );
  AOI221_X1 U2009 ( .B1(n6240), .B2(\registers[13][17] ), .C1(n6244), .C2(
        \registers[12][17] ), .A(n5400), .ZN(n5397) );
  OAI22_X1 U2010 ( .A1(n2828), .A2(n6249), .B1(n5818), .B2(n6257), .ZN(n5400)
         );
  AOI221_X1 U2011 ( .B1(n5116), .B2(\registers[31][17] ), .C1(n5117), .C2(
        \registers[30][17] ), .A(n5402), .ZN(n5395) );
  OAI22_X1 U2012 ( .A1(n4174), .A2(n6191), .B1(n5876), .B2(n6198), .ZN(n5402)
         );
  AOI221_X1 U2013 ( .B1(n6208), .B2(\registers[21][17] ), .C1(n6216), .C2(
        \registers[20][17] ), .A(n5401), .ZN(n5396) );
  OAI22_X1 U2014 ( .A1(n2829), .A2(n6221), .B1(n5819), .B2(n6231), .ZN(n5401)
         );
  AOI221_X1 U2015 ( .B1(n6114), .B2(\registers[29][17] ), .C1(n6118), .C2(
        \registers[28][17] ), .A(n5409), .ZN(n5404) );
  OAI22_X1 U2016 ( .A1(n4237), .A2(n6121), .B1(n5935), .B2(n6130), .ZN(n5409)
         );
  AOI221_X1 U2017 ( .B1(n6082), .B2(\registers[23][17] ), .C1(n6090), .C2(
        \registers[22][17] ), .A(n5410), .ZN(n5403) );
  OAI22_X1 U2018 ( .A1(n4175), .A2(n6096), .B1(n5877), .B2(n6104), .ZN(n5410)
         );
  AOI221_X1 U2019 ( .B1(n6241), .B2(\registers[13][18] ), .C1(n6243), .C2(
        \registers[12][18] ), .A(n5381), .ZN(n5378) );
  OAI22_X1 U2020 ( .A1(n2830), .A2(n6250), .B1(n5820), .B2(n6258), .ZN(n5381)
         );
  AOI221_X1 U2021 ( .B1(n6182), .B2(\registers[31][18] ), .C1(n6184), .C2(
        \registers[30][18] ), .A(n5383), .ZN(n5376) );
  OAI22_X1 U2022 ( .A1(n4176), .A2(n6192), .B1(n5878), .B2(n6199), .ZN(n5383)
         );
  AOI221_X1 U2023 ( .B1(n6209), .B2(\registers[21][18] ), .C1(n6216), .C2(
        \registers[20][18] ), .A(n5382), .ZN(n5377) );
  OAI22_X1 U2024 ( .A1(n2831), .A2(n6224), .B1(n5821), .B2(n6228), .ZN(n5382)
         );
  AOI221_X1 U2025 ( .B1(n6115), .B2(\registers[29][18] ), .C1(n6117), .C2(
        \registers[28][18] ), .A(n5390), .ZN(n5385) );
  OAI22_X1 U2026 ( .A1(n4238), .A2(n6124), .B1(n5936), .B2(n6132), .ZN(n5390)
         );
  AOI221_X1 U2027 ( .B1(n6083), .B2(\registers[23][18] ), .C1(n6091), .C2(
        \registers[22][18] ), .A(n5391), .ZN(n5384) );
  OAI22_X1 U2028 ( .A1(n4177), .A2(n6097), .B1(n5879), .B2(n6106), .ZN(n5391)
         );
  AOI221_X1 U2029 ( .B1(n6241), .B2(\registers[13][19] ), .C1(n6244), .C2(
        \registers[12][19] ), .A(n5362), .ZN(n5359) );
  OAI22_X1 U2030 ( .A1(n2832), .A2(n6251), .B1(n5822), .B2(n6260), .ZN(n5362)
         );
  AOI221_X1 U2031 ( .B1(n6183), .B2(\registers[31][19] ), .C1(n6185), .C2(
        \registers[30][19] ), .A(n5364), .ZN(n5357) );
  OAI22_X1 U2032 ( .A1(n4178), .A2(n6193), .B1(n5880), .B2(n6200), .ZN(n5364)
         );
  AOI221_X1 U2033 ( .B1(n6209), .B2(\registers[21][19] ), .C1(n6217), .C2(
        \registers[20][19] ), .A(n5363), .ZN(n5358) );
  OAI22_X1 U2034 ( .A1(n2833), .A2(n6225), .B1(n5823), .B2(n6232), .ZN(n5363)
         );
  AOI221_X1 U2035 ( .B1(n6115), .B2(\registers[29][19] ), .C1(n6118), .C2(
        \registers[28][19] ), .A(n5371), .ZN(n5366) );
  OAI22_X1 U2036 ( .A1(n4239), .A2(n6125), .B1(n5937), .B2(n6133), .ZN(n5371)
         );
  AOI221_X1 U2037 ( .B1(n6083), .B2(\registers[23][19] ), .C1(n6091), .C2(
        \registers[22][19] ), .A(n5372), .ZN(n5365) );
  OAI22_X1 U2038 ( .A1(n4179), .A2(n6098), .B1(n5881), .B2(n6105), .ZN(n5372)
         );
  AOI221_X1 U2039 ( .B1(n6241), .B2(\registers[13][20] ), .C1(n6242), .C2(
        \registers[12][20] ), .A(n5343), .ZN(n5340) );
  OAI22_X1 U2040 ( .A1(n2834), .A2(n6250), .B1(n5824), .B2(n6259), .ZN(n5343)
         );
  AOI221_X1 U2041 ( .B1(n6209), .B2(\registers[21][20] ), .C1(n6217), .C2(
        \registers[20][20] ), .A(n5344), .ZN(n5339) );
  OAI22_X1 U2042 ( .A1(n2835), .A2(n6220), .B1(n5825), .B2(n6233), .ZN(n5344)
         );
  AOI221_X1 U2043 ( .B1(n6115), .B2(\registers[29][20] ), .C1(n6116), .C2(
        \registers[28][20] ), .A(n5352), .ZN(n5347) );
  OAI22_X1 U2044 ( .A1(n4240), .A2(n6125), .B1(n5938), .B2(n6134), .ZN(n5352)
         );
  AOI221_X1 U2045 ( .B1(n6083), .B2(\registers[23][20] ), .C1(n6091), .C2(
        \registers[22][20] ), .A(n5353), .ZN(n5346) );
  OAI22_X1 U2046 ( .A1(n4180), .A2(n6099), .B1(n5882), .B2(n6105), .ZN(n5353)
         );
  AOI221_X1 U2047 ( .B1(n6241), .B2(\registers[13][21] ), .C1(n6242), .C2(
        \registers[12][21] ), .A(n5324), .ZN(n5321) );
  OAI22_X1 U2048 ( .A1(n2836), .A2(n6252), .B1(n5826), .B2(n6260), .ZN(n5324)
         );
  AOI221_X1 U2049 ( .B1(n6209), .B2(\registers[21][21] ), .C1(n6217), .C2(
        \registers[20][21] ), .A(n5325), .ZN(n5320) );
  OAI22_X1 U2050 ( .A1(n2837), .A2(n6224), .B1(n5827), .B2(n6233), .ZN(n5325)
         );
  AOI221_X1 U2051 ( .B1(n6115), .B2(\registers[29][21] ), .C1(n6116), .C2(
        \registers[28][21] ), .A(n5333), .ZN(n5328) );
  OAI22_X1 U2052 ( .A1(n4241), .A2(n6126), .B1(n5939), .B2(n6134), .ZN(n5333)
         );
  AOI221_X1 U2053 ( .B1(n6083), .B2(\registers[23][21] ), .C1(n6091), .C2(
        \registers[22][21] ), .A(n5334), .ZN(n5327) );
  OAI22_X1 U2054 ( .A1(n4181), .A2(n6097), .B1(n5883), .B2(n6105), .ZN(n5334)
         );
  AOI221_X1 U2055 ( .B1(n6235), .B2(\registers[13][22] ), .C1(n6243), .C2(
        \registers[12][22] ), .A(n5305), .ZN(n5302) );
  OAI22_X1 U2056 ( .A1(n2838), .A2(n6252), .B1(n5828), .B2(n6258), .ZN(n5305)
         );
  AOI221_X1 U2057 ( .B1(n6077), .B2(\registers[23][22] ), .C1(n6086), .C2(
        \registers[22][22] ), .A(n5315), .ZN(n5308) );
  OAI22_X1 U2058 ( .A1(n4185), .A2(n6099), .B1(n5884), .B2(n6106), .ZN(n5315)
         );
  AOI221_X1 U2059 ( .B1(n6236), .B2(\registers[13][23] ), .C1(n6243), .C2(
        \registers[12][23] ), .A(n5286), .ZN(n5283) );
  OAI22_X1 U2060 ( .A1(n2839), .A2(n6251), .B1(n5829), .B2(n6259), .ZN(n5286)
         );
  AOI221_X1 U2061 ( .B1(n6078), .B2(\registers[23][23] ), .C1(n6085), .C2(
        \registers[22][23] ), .A(n5296), .ZN(n5289) );
  OAI22_X1 U2062 ( .A1(n4186), .A2(n6093), .B1(n5885), .B2(n6107), .ZN(n5296)
         );
  AOI221_X1 U2063 ( .B1(n6235), .B2(\registers[13][24] ), .C1(n6244), .C2(
        \registers[12][24] ), .A(n5267), .ZN(n5264) );
  OAI22_X1 U2064 ( .A1(n2840), .A2(n6246), .B1(n5830), .B2(n6255), .ZN(n5267)
         );
  AOI221_X1 U2065 ( .B1(n6078), .B2(\registers[23][24] ), .C1(n6085), .C2(
        \registers[22][24] ), .A(n5277), .ZN(n5270) );
  OAI22_X1 U2066 ( .A1(n4187), .A2(n6097), .B1(n5886), .B2(n6103), .ZN(n5277)
         );
  AOI221_X1 U2067 ( .B1(n6237), .B2(\registers[13][25] ), .C1(n6242), .C2(
        \registers[12][25] ), .A(n5248), .ZN(n5245) );
  OAI22_X1 U2068 ( .A1(n2841), .A2(n6246), .B1(n5831), .B2(n6260), .ZN(n5248)
         );
  AOI221_X1 U2069 ( .B1(n6079), .B2(\registers[23][25] ), .C1(n6086), .C2(
        \registers[22][25] ), .A(n5258), .ZN(n5251) );
  OAI22_X1 U2070 ( .A1(n4188), .A2(n6099), .B1(n5887), .B2(n6107), .ZN(n5258)
         );
  AOI221_X1 U2071 ( .B1(n6237), .B2(\registers[13][26] ), .C1(n6244), .C2(
        \registers[12][26] ), .A(n5229), .ZN(n5226) );
  OAI22_X1 U2072 ( .A1(n2842), .A2(n6252), .B1(n5832), .B2(n6256), .ZN(n5229)
         );
  AOI221_X1 U2073 ( .B1(n6079), .B2(\registers[23][26] ), .C1(n6086), .C2(
        \registers[22][26] ), .A(n5239), .ZN(n5232) );
  OAI22_X1 U2074 ( .A1(n4189), .A2(n6098), .B1(n5888), .B2(n6102), .ZN(n5239)
         );
  AOI221_X1 U2075 ( .B1(n6235), .B2(\registers[13][27] ), .C1(n6243), .C2(
        \registers[12][27] ), .A(n5210), .ZN(n5207) );
  OAI22_X1 U2076 ( .A1(n2843), .A2(n6252), .B1(n5833), .B2(n6260), .ZN(n5210)
         );
  AOI221_X1 U2077 ( .B1(n6077), .B2(\registers[23][27] ), .C1(n6089), .C2(
        \registers[22][27] ), .A(n5220), .ZN(n5213) );
  OAI22_X1 U2078 ( .A1(n4190), .A2(n6098), .B1(n5889), .B2(n6106), .ZN(n5220)
         );
  AOI221_X1 U2079 ( .B1(n6238), .B2(\registers[13][28] ), .C1(n6244), .C2(
        \registers[12][28] ), .A(n5191), .ZN(n5188) );
  OAI22_X1 U2080 ( .A1(n2844), .A2(n6248), .B1(n5834), .B2(n6254), .ZN(n5191)
         );
  AOI221_X1 U2081 ( .B1(n6183), .B2(\registers[31][28] ), .C1(n6185), .C2(
        \registers[30][28] ), .A(n5193), .ZN(n5186) );
  OAI22_X1 U2082 ( .A1(n4191), .A2(n6187), .B1(n5890), .B2(n6201), .ZN(n5193)
         );
  AOI221_X1 U2083 ( .B1(n6205), .B2(\registers[21][28] ), .C1(n6213), .C2(
        \registers[20][28] ), .A(n5192), .ZN(n5187) );
  OAI22_X1 U2084 ( .A1(n2845), .A2(n6219), .B1(n5835), .B2(n6227), .ZN(n5192)
         );
  AOI221_X1 U2085 ( .B1(n6110), .B2(\registers[29][28] ), .C1(n6118), .C2(
        \registers[28][28] ), .A(n5200), .ZN(n5195) );
  OAI22_X1 U2086 ( .A1(n4242), .A2(n6126), .B1(n5940), .B2(n6128), .ZN(n5200)
         );
  AOI221_X1 U2087 ( .B1(n6080), .B2(\registers[23][28] ), .C1(n6085), .C2(
        \registers[22][28] ), .A(n5201), .ZN(n5194) );
  OAI22_X1 U2088 ( .A1(n4192), .A2(n6095), .B1(n5891), .B2(n6101), .ZN(n5201)
         );
  AOI221_X1 U2089 ( .B1(n6236), .B2(\registers[13][29] ), .C1(n6242), .C2(
        \registers[12][29] ), .A(n5172), .ZN(n5169) );
  OAI22_X1 U2090 ( .A1(n2846), .A2(n6252), .B1(n5836), .B2(n6258), .ZN(n5172)
         );
  AOI221_X1 U2091 ( .B1(n5116), .B2(\registers[31][29] ), .C1(n5117), .C2(
        \registers[30][29] ), .A(n5174), .ZN(n5167) );
  OAI22_X1 U2092 ( .A1(n4193), .A2(n6189), .B1(n5892), .B2(n6196), .ZN(n5174)
         );
  AOI221_X1 U2093 ( .B1(n6204), .B2(\registers[21][29] ), .C1(n6213), .C2(
        \registers[20][29] ), .A(n5173), .ZN(n5168) );
  OAI22_X1 U2094 ( .A1(n2847), .A2(n6223), .B1(n5837), .B2(n6231), .ZN(n5173)
         );
  AOI221_X1 U2095 ( .B1(n6111), .B2(\registers[29][29] ), .C1(n6116), .C2(
        \registers[28][29] ), .A(n5181), .ZN(n5176) );
  OAI22_X1 U2096 ( .A1(n4243), .A2(n6123), .B1(n5941), .B2(n6131), .ZN(n5181)
         );
  AOI221_X1 U2097 ( .B1(n6078), .B2(\registers[23][29] ), .C1(n6087), .C2(
        \registers[22][29] ), .A(n5182), .ZN(n5175) );
  OAI22_X1 U2098 ( .A1(n4194), .A2(n6099), .B1(n5893), .B2(n6106), .ZN(n5182)
         );
  AOI221_X1 U2099 ( .B1(n6236), .B2(\registers[13][30] ), .C1(n6242), .C2(
        \registers[12][30] ), .A(n5153), .ZN(n5150) );
  OAI22_X1 U2100 ( .A1(n2848), .A2(n6250), .B1(n5838), .B2(n6254), .ZN(n5153)
         );
  AOI221_X1 U2101 ( .B1(n6182), .B2(\registers[31][30] ), .C1(n6184), .C2(
        \registers[30][30] ), .A(n5155), .ZN(n5148) );
  OAI22_X1 U2102 ( .A1(n4195), .A2(n6188), .B1(n5894), .B2(n6200), .ZN(n5155)
         );
  AOI221_X1 U2103 ( .B1(n6203), .B2(\registers[21][30] ), .C1(n6214), .C2(
        \registers[20][30] ), .A(n5154), .ZN(n5149) );
  OAI22_X1 U2104 ( .A1(n2849), .A2(n6225), .B1(n5839), .B2(n6228), .ZN(n5154)
         );
  AOI221_X1 U2105 ( .B1(n6111), .B2(\registers[29][30] ), .C1(n6116), .C2(
        \registers[28][30] ), .A(n5162), .ZN(n5157) );
  OAI22_X1 U2106 ( .A1(n4244), .A2(n6120), .B1(n5942), .B2(n6133), .ZN(n5162)
         );
  AOI221_X1 U2107 ( .B1(n6078), .B2(\registers[23][30] ), .C1(n6087), .C2(
        \registers[22][30] ), .A(n5163), .ZN(n5156) );
  OAI22_X1 U2108 ( .A1(n4196), .A2(n6099), .B1(n5895), .B2(n6105), .ZN(n5163)
         );
  AOI221_X1 U2109 ( .B1(n6238), .B2(\registers[13][31] ), .C1(n6243), .C2(
        \registers[12][31] ), .A(n5108), .ZN(n5099) );
  OAI22_X1 U2110 ( .A1(n2850), .A2(n6246), .B1(n5840), .B2(n6254), .ZN(n5108)
         );
  AOI221_X1 U2111 ( .B1(n6183), .B2(\registers[31][31] ), .C1(n6185), .C2(
        \registers[30][31] ), .A(n5118), .ZN(n5097) );
  OAI22_X1 U2112 ( .A1(n4197), .A2(n6192), .B1(n5896), .B2(n6195), .ZN(n5118)
         );
  AOI221_X1 U2113 ( .B1(n6206), .B2(\registers[21][31] ), .C1(n6213), .C2(
        \registers[20][31] ), .A(n5113), .ZN(n5098) );
  OAI22_X1 U2114 ( .A1(n2851), .A2(n6224), .B1(n5841), .B2(n6233), .ZN(n5113)
         );
  AOI221_X1 U2115 ( .B1(n6112), .B2(\registers[29][31] ), .C1(n6117), .C2(
        \registers[28][31] ), .A(n5137), .ZN(n5122) );
  OAI22_X1 U2116 ( .A1(n4245), .A2(n6125), .B1(n5943), .B2(n6128), .ZN(n5137)
         );
  AOI221_X1 U2117 ( .B1(n6080), .B2(\registers[23][31] ), .C1(n6088), .C2(
        \registers[22][31] ), .A(n5142), .ZN(n5121) );
  OAI22_X1 U2118 ( .A1(n4198), .A2(n6097), .B1(n5897), .B2(n6107), .ZN(n5142)
         );
  AOI221_X1 U2119 ( .B1(\registers[31][0] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][0] ), .A(n5066), .ZN(n5051) );
  OAI22_X1 U2120 ( .A1(n2852), .A2(n6400), .B1(n5842), .B2(n6406), .ZN(n5066)
         );
  AOI221_X1 U2121 ( .B1(n6282), .B2(\registers[23][0] ), .C1(n6290), .C2(
        \registers[22][0] ), .A(n5082), .ZN(n5071) );
  OAI22_X1 U2122 ( .A1(n2853), .A2(n6294), .B1(n5843), .B2(n6307), .ZN(n5082)
         );
  AOI221_X1 U2123 ( .B1(n6309), .B2(\registers[25][0] ), .C1(n6320), .C2(
        \registers[24][0] ), .A(n5079), .ZN(n5072) );
  OAI22_X1 U2124 ( .A1(n4246), .A2(n6325), .B1(n5944), .B2(n6333), .ZN(n5079)
         );
  AOI221_X1 U2125 ( .B1(\registers[31][1] ), .B2(n6392), .C1(n6394), .C2(
        \registers[30][1] ), .A(n5037), .ZN(n5030) );
  OAI22_X1 U2126 ( .A1(n2854), .A2(n6402), .B1(n5844), .B2(n6404), .ZN(n5037)
         );
  AOI221_X1 U2127 ( .B1(n6283), .B2(\registers[23][1] ), .C1(n6291), .C2(
        \registers[22][1] ), .A(n5045), .ZN(n5038) );
  OAI22_X1 U2128 ( .A1(n2855), .A2(n6297), .B1(n5845), .B2(n6307), .ZN(n5045)
         );
  AOI221_X1 U2129 ( .B1(n6310), .B2(\registers[25][1] ), .C1(n6320), .C2(
        \registers[24][1] ), .A(n5044), .ZN(n5039) );
  OAI22_X1 U2130 ( .A1(n4247), .A2(n6327), .B1(n5945), .B2(n6334), .ZN(n5044)
         );
  AOI221_X1 U2131 ( .B1(\registers[31][2] ), .B2(n4417), .C1(n4418), .C2(
        \registers[30][2] ), .A(n5017), .ZN(n5010) );
  OAI22_X1 U2132 ( .A1(n2856), .A2(n6398), .B1(n5846), .B2(n6407), .ZN(n5017)
         );
  AOI221_X1 U2133 ( .B1(n6282), .B2(\registers[23][2] ), .C1(n6289), .C2(
        \registers[22][2] ), .A(n5025), .ZN(n5018) );
  OAI22_X1 U2134 ( .A1(n2857), .A2(n6299), .B1(n5847), .B2(n6305), .ZN(n5025)
         );
  AOI221_X1 U2135 ( .B1(n6309), .B2(\registers[25][2] ), .C1(n6317), .C2(
        \registers[24][2] ), .A(n5024), .ZN(n5019) );
  OAI22_X1 U2136 ( .A1(n4248), .A2(n6329), .B1(n5946), .B2(n6333), .ZN(n5024)
         );
  AOI221_X1 U2137 ( .B1(\registers[31][3] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][3] ), .A(n4997), .ZN(n4990) );
  OAI22_X1 U2138 ( .A1(n2860), .A2(n6397), .B1(n5848), .B2(n6408), .ZN(n4997)
         );
  AOI221_X1 U2139 ( .B1(n6284), .B2(\registers[23][3] ), .C1(n6289), .C2(
        \registers[22][3] ), .A(n5005), .ZN(n4998) );
  OAI22_X1 U2140 ( .A1(n2895), .A2(n6297), .B1(n5849), .B2(n6305), .ZN(n5005)
         );
  AOI221_X1 U2141 ( .B1(n6311), .B2(\registers[25][3] ), .C1(n6318), .C2(
        \registers[24][3] ), .A(n5004), .ZN(n4999) );
  OAI22_X1 U2142 ( .A1(n4249), .A2(n6326), .B1(n5947), .B2(n6334), .ZN(n5004)
         );
  AOI221_X1 U2143 ( .B1(\registers[31][4] ), .B2(n6392), .C1(n6394), .C2(
        \registers[30][4] ), .A(n4977), .ZN(n4970) );
  OAI22_X1 U2144 ( .A1(n2929), .A2(n6396), .B1(n5850), .B2(n6404), .ZN(n4977)
         );
  AOI221_X1 U2145 ( .B1(n6285), .B2(\registers[23][4] ), .C1(n6290), .C2(
        \registers[22][4] ), .A(n4985), .ZN(n4978) );
  OAI22_X1 U2146 ( .A1(n2971), .A2(n6293), .B1(n5851), .B2(n6301), .ZN(n4985)
         );
  AOI221_X1 U2147 ( .B1(n6312), .B2(\registers[25][4] ), .C1(n6318), .C2(
        \registers[24][4] ), .A(n4984), .ZN(n4979) );
  OAI22_X1 U2148 ( .A1(n4250), .A2(n6326), .B1(n5948), .B2(n6335), .ZN(n4984)
         );
  AOI221_X1 U2149 ( .B1(\registers[31][5] ), .B2(n4417), .C1(n4418), .C2(
        \registers[30][5] ), .A(n4957), .ZN(n4950) );
  OAI22_X1 U2150 ( .A1(n4150), .A2(n6397), .B1(n5852), .B2(n6405), .ZN(n4957)
         );
  AOI221_X1 U2151 ( .B1(n6284), .B2(\registers[23][5] ), .C1(n6290), .C2(
        \registers[22][5] ), .A(n4965), .ZN(n4958) );
  OAI22_X1 U2152 ( .A1(n4151), .A2(n6294), .B1(n5853), .B2(n6302), .ZN(n4965)
         );
  AOI221_X1 U2153 ( .B1(n6311), .B2(\registers[25][5] ), .C1(n6322), .C2(
        \registers[24][5] ), .A(n4964), .ZN(n4959) );
  OAI22_X1 U2154 ( .A1(n4253), .A2(n6326), .B1(n5949), .B2(n6336), .ZN(n4964)
         );
  AOI221_X1 U2155 ( .B1(\registers[31][6] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][6] ), .A(n4937), .ZN(n4930) );
  OAI22_X1 U2156 ( .A1(n4152), .A2(n6398), .B1(n5854), .B2(n6406), .ZN(n4937)
         );
  AOI221_X1 U2157 ( .B1(n6288), .B2(\registers[23][6] ), .C1(n6291), .C2(
        \registers[22][6] ), .A(n4945), .ZN(n4938) );
  OAI22_X1 U2158 ( .A1(n4153), .A2(n6295), .B1(n5855), .B2(n6303), .ZN(n4945)
         );
  AOI221_X1 U2159 ( .B1(n6315), .B2(\registers[25][6] ), .C1(n6319), .C2(
        \registers[24][6] ), .A(n4944), .ZN(n4939) );
  OAI22_X1 U2160 ( .A1(n4254), .A2(n6327), .B1(n5950), .B2(n6335), .ZN(n4944)
         );
  AOI221_X1 U2161 ( .B1(\registers[31][7] ), .B2(n6392), .C1(n6394), .C2(
        \registers[30][7] ), .A(n4917), .ZN(n4910) );
  OAI22_X1 U2162 ( .A1(n4154), .A2(n6399), .B1(n5856), .B2(n6407), .ZN(n4917)
         );
  AOI221_X1 U2163 ( .B1(n6286), .B2(\registers[23][7] ), .C1(n6289), .C2(
        \registers[22][7] ), .A(n4925), .ZN(n4918) );
  OAI22_X1 U2164 ( .A1(n4155), .A2(n6296), .B1(n5857), .B2(n6304), .ZN(n4925)
         );
  AOI221_X1 U2165 ( .B1(n6313), .B2(\registers[25][7] ), .C1(n6319), .C2(
        \registers[24][7] ), .A(n4924), .ZN(n4919) );
  OAI22_X1 U2166 ( .A1(n4255), .A2(n6328), .B1(n5951), .B2(n6336), .ZN(n4924)
         );
  AOI221_X1 U2167 ( .B1(\registers[31][8] ), .B2(n4417), .C1(n4418), .C2(
        \registers[30][8] ), .A(n4897), .ZN(n4890) );
  OAI22_X1 U2168 ( .A1(n4156), .A2(n6400), .B1(n5858), .B2(n6408), .ZN(n4897)
         );
  AOI221_X1 U2169 ( .B1(n6286), .B2(\registers[23][8] ), .C1(n6291), .C2(
        \registers[22][8] ), .A(n4905), .ZN(n4898) );
  OAI22_X1 U2170 ( .A1(n4157), .A2(n6296), .B1(n5859), .B2(n6302), .ZN(n4905)
         );
  AOI221_X1 U2171 ( .B1(n6313), .B2(\registers[25][8] ), .C1(n6321), .C2(
        \registers[24][8] ), .A(n4904), .ZN(n4899) );
  OAI22_X1 U2172 ( .A1(n4256), .A2(n6328), .B1(n5952), .B2(n6337), .ZN(n4904)
         );
  AOI221_X1 U2173 ( .B1(\registers[31][9] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][9] ), .A(n4877), .ZN(n4870) );
  OAI22_X1 U2174 ( .A1(n4158), .A2(n6401), .B1(n5860), .B2(n6409), .ZN(n4877)
         );
  AOI221_X1 U2175 ( .B1(n6286), .B2(\registers[23][9] ), .C1(n6290), .C2(
        \registers[22][9] ), .A(n4885), .ZN(n4878) );
  OAI22_X1 U2176 ( .A1(n4159), .A2(n6296), .B1(n5861), .B2(n6304), .ZN(n4885)
         );
  AOI221_X1 U2177 ( .B1(n6313), .B2(\registers[25][9] ), .C1(n6321), .C2(
        \registers[24][9] ), .A(n4884), .ZN(n4879) );
  OAI22_X1 U2178 ( .A1(n4257), .A2(n6327), .B1(n5953), .B2(n6338), .ZN(n4884)
         );
  AOI221_X1 U2179 ( .B1(\registers[31][10] ), .B2(n6392), .C1(n6394), .C2(
        \registers[30][10] ), .A(n4857), .ZN(n4850) );
  OAI22_X1 U2180 ( .A1(n4160), .A2(n6398), .B1(n5862), .B2(n6408), .ZN(n4857)
         );
  AOI221_X1 U2181 ( .B1(n6285), .B2(\registers[23][10] ), .C1(n6291), .C2(
        \registers[22][10] ), .A(n4865), .ZN(n4858) );
  OAI22_X1 U2182 ( .A1(n4161), .A2(n6297), .B1(n5863), .B2(n6305), .ZN(n4865)
         );
  AOI221_X1 U2183 ( .B1(n6312), .B2(\registers[25][10] ), .C1(n6320), .C2(
        \registers[24][10] ), .A(n4864), .ZN(n4859) );
  OAI22_X1 U2184 ( .A1(n4258), .A2(n6329), .B1(n5954), .B2(n6333), .ZN(n4864)
         );
  AOI221_X1 U2185 ( .B1(\registers[31][11] ), .B2(n4417), .C1(n4418), .C2(
        \registers[30][11] ), .A(n4837), .ZN(n4830) );
  OAI22_X1 U2186 ( .A1(n4162), .A2(n6396), .B1(n5864), .B2(n6404), .ZN(n4837)
         );
  AOI221_X1 U2187 ( .B1(n6286), .B2(\registers[23][11] ), .C1(n6289), .C2(
        \registers[22][11] ), .A(n4845), .ZN(n4838) );
  OAI22_X1 U2188 ( .A1(n4163), .A2(n6298), .B1(n5865), .B2(n6301), .ZN(n4845)
         );
  AOI221_X1 U2189 ( .B1(n6313), .B2(\registers[25][11] ), .C1(n6321), .C2(
        \registers[24][11] ), .A(n4844), .ZN(n4839) );
  OAI22_X1 U2190 ( .A1(n4259), .A2(n6330), .B1(n5955), .B2(n6334), .ZN(n4844)
         );
  AOI221_X1 U2191 ( .B1(\registers[31][12] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][12] ), .A(n4817), .ZN(n4810) );
  OAI22_X1 U2192 ( .A1(n4164), .A2(n6396), .B1(n5866), .B2(n6404), .ZN(n4817)
         );
  AOI221_X1 U2193 ( .B1(n6287), .B2(\registers[23][12] ), .C1(n6289), .C2(
        \registers[22][12] ), .A(n4825), .ZN(n4818) );
  OAI22_X1 U2194 ( .A1(n4165), .A2(n6293), .B1(n5867), .B2(n6301), .ZN(n4825)
         );
  AOI221_X1 U2195 ( .B1(n6314), .B2(\registers[25][12] ), .C1(n6322), .C2(
        \registers[24][12] ), .A(n4824), .ZN(n4819) );
  OAI22_X1 U2196 ( .A1(n4260), .A2(n6326), .B1(n5956), .B2(n6337), .ZN(n4824)
         );
  AOI221_X1 U2197 ( .B1(\registers[31][13] ), .B2(n6392), .C1(n6394), .C2(
        \registers[30][13] ), .A(n4797), .ZN(n4790) );
  OAI22_X1 U2198 ( .A1(n4166), .A2(n6397), .B1(n5868), .B2(n6405), .ZN(n4797)
         );
  AOI221_X1 U2199 ( .B1(n6287), .B2(\registers[23][13] ), .C1(n6290), .C2(
        \registers[22][13] ), .A(n4805), .ZN(n4798) );
  OAI22_X1 U2200 ( .A1(n4167), .A2(n6294), .B1(n5869), .B2(n6302), .ZN(n4805)
         );
  AOI221_X1 U2201 ( .B1(n6314), .B2(\registers[25][13] ), .C1(n6322), .C2(
        \registers[24][13] ), .A(n4804), .ZN(n4799) );
  OAI22_X1 U2202 ( .A1(n4261), .A2(n6326), .B1(n5957), .B2(n6338), .ZN(n4804)
         );
  AOI221_X1 U2203 ( .B1(\registers[31][14] ), .B2(n4417), .C1(n4418), .C2(
        \registers[30][14] ), .A(n4777), .ZN(n4770) );
  OAI22_X1 U2204 ( .A1(n4168), .A2(n6398), .B1(n5870), .B2(n6406), .ZN(n4777)
         );
  AOI221_X1 U2205 ( .B1(n6285), .B2(\registers[23][14] ), .C1(n6290), .C2(
        \registers[22][14] ), .A(n4785), .ZN(n4778) );
  OAI22_X1 U2206 ( .A1(n4169), .A2(n6295), .B1(n5871), .B2(n6303), .ZN(n4785)
         );
  AOI221_X1 U2207 ( .B1(n6312), .B2(\registers[25][14] ), .C1(n6320), .C2(
        \registers[24][14] ), .A(n4784), .ZN(n4779) );
  OAI22_X1 U2208 ( .A1(n4262), .A2(n6327), .B1(n5958), .B2(n6335), .ZN(n4784)
         );
  AOI221_X1 U2209 ( .B1(\registers[31][15] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][15] ), .A(n4757), .ZN(n4750) );
  OAI22_X1 U2210 ( .A1(n4170), .A2(n6399), .B1(n5872), .B2(n6407), .ZN(n4757)
         );
  AOI221_X1 U2211 ( .B1(n6286), .B2(\registers[23][15] ), .C1(n6291), .C2(
        \registers[22][15] ), .A(n4765), .ZN(n4758) );
  OAI22_X1 U2212 ( .A1(n4171), .A2(n6296), .B1(n5873), .B2(n6303), .ZN(n4765)
         );
  AOI221_X1 U2213 ( .B1(n6313), .B2(\registers[25][15] ), .C1(n6321), .C2(
        \registers[24][15] ), .A(n4764), .ZN(n4759) );
  OAI22_X1 U2214 ( .A1(n4263), .A2(n6328), .B1(n5959), .B2(n6336), .ZN(n4764)
         );
  AOI221_X1 U2215 ( .B1(\registers[31][16] ), .B2(n6392), .C1(n6394), .C2(
        \registers[30][16] ), .A(n4737), .ZN(n4730) );
  OAI22_X1 U2216 ( .A1(n4172), .A2(n6400), .B1(n5874), .B2(n6408), .ZN(n4737)
         );
  AOI221_X1 U2217 ( .B1(n6287), .B2(\registers[23][16] ), .C1(n6289), .C2(
        \registers[22][16] ), .A(n4745), .ZN(n4738) );
  OAI22_X1 U2218 ( .A1(n4173), .A2(n6295), .B1(n5875), .B2(n6303), .ZN(n4745)
         );
  AOI221_X1 U2219 ( .B1(n6314), .B2(\registers[25][16] ), .C1(n6322), .C2(
        \registers[24][16] ), .A(n4744), .ZN(n4739) );
  OAI22_X1 U2220 ( .A1(n4264), .A2(n6328), .B1(n5960), .B2(n6337), .ZN(n4744)
         );
  AOI221_X1 U2221 ( .B1(\registers[31][17] ), .B2(n4417), .C1(n4418), .C2(
        \registers[30][17] ), .A(n4717), .ZN(n4710) );
  OAI22_X1 U2222 ( .A1(n4174), .A2(n6401), .B1(n5876), .B2(n6409), .ZN(n4717)
         );
  AOI221_X1 U2223 ( .B1(n6287), .B2(\registers[23][17] ), .C1(n6291), .C2(
        \registers[22][17] ), .A(n4725), .ZN(n4718) );
  OAI22_X1 U2224 ( .A1(n4175), .A2(n6294), .B1(n5877), .B2(n6304), .ZN(n4725)
         );
  AOI221_X1 U2225 ( .B1(n6314), .B2(\registers[25][17] ), .C1(n6322), .C2(
        \registers[24][17] ), .A(n4724), .ZN(n4719) );
  OAI22_X1 U2226 ( .A1(n4265), .A2(n6327), .B1(n5961), .B2(n6338), .ZN(n4724)
         );
  AOI221_X1 U2227 ( .B1(\registers[31][18] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][18] ), .A(n4697), .ZN(n4690) );
  OAI22_X1 U2228 ( .A1(n4176), .A2(n6396), .B1(n5878), .B2(n6408), .ZN(n4697)
         );
  AOI221_X1 U2229 ( .B1(n6288), .B2(\registers[23][18] ), .C1(n6290), .C2(
        \registers[22][18] ), .A(n4705), .ZN(n4698) );
  OAI22_X1 U2230 ( .A1(n4177), .A2(n6297), .B1(n5879), .B2(n6305), .ZN(n4705)
         );
  AOI221_X1 U2231 ( .B1(n6315), .B2(\registers[25][18] ), .C1(n6323), .C2(
        \registers[24][18] ), .A(n4704), .ZN(n4699) );
  OAI22_X1 U2232 ( .A1(n4266), .A2(n6329), .B1(n5962), .B2(n6333), .ZN(n4704)
         );
  AOI221_X1 U2233 ( .B1(\registers[31][19] ), .B2(n6392), .C1(n6394), .C2(
        \registers[30][19] ), .A(n4677), .ZN(n4670) );
  OAI22_X1 U2234 ( .A1(n4178), .A2(n6400), .B1(n5880), .B2(n6406), .ZN(n4677)
         );
  AOI221_X1 U2235 ( .B1(n6288), .B2(\registers[23][19] ), .C1(n6291), .C2(
        \registers[22][19] ), .A(n4685), .ZN(n4678) );
  OAI22_X1 U2236 ( .A1(n4179), .A2(n6298), .B1(n5881), .B2(n6307), .ZN(n4685)
         );
  AOI221_X1 U2237 ( .B1(n6315), .B2(\registers[25][19] ), .C1(n6323), .C2(
        \registers[24][19] ), .A(n4684), .ZN(n4679) );
  OAI22_X1 U2238 ( .A1(n4267), .A2(n6330), .B1(n5963), .B2(n6334), .ZN(n4684)
         );
  AOI221_X1 U2239 ( .B1(\registers[31][20] ), .B2(n4417), .C1(n4418), .C2(
        \registers[30][20] ), .A(n4657), .ZN(n4650) );
  OAI22_X1 U2240 ( .A1(n4199), .A2(n6396), .B1(n5898), .B2(n6410), .ZN(n4657)
         );
  AOI221_X1 U2241 ( .B1(n6288), .B2(\registers[23][20] ), .C1(n6289), .C2(
        \registers[22][20] ), .A(n4665), .ZN(n4658) );
  OAI22_X1 U2242 ( .A1(n4180), .A2(n6298), .B1(n5882), .B2(n6306), .ZN(n4665)
         );
  AOI221_X1 U2243 ( .B1(n6315), .B2(\registers[25][20] ), .C1(n6323), .C2(
        \registers[24][20] ), .A(n4664), .ZN(n4659) );
  OAI22_X1 U2244 ( .A1(n4268), .A2(n6331), .B1(n5964), .B2(n6333), .ZN(n4664)
         );
  AOI221_X1 U2245 ( .B1(\registers[31][21] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][21] ), .A(n4637), .ZN(n4630) );
  OAI22_X1 U2246 ( .A1(n4200), .A2(n6402), .B1(n5899), .B2(n6410), .ZN(n4637)
         );
  AOI221_X1 U2247 ( .B1(n6288), .B2(\registers[23][21] ), .C1(n6289), .C2(
        \registers[22][21] ), .A(n4645), .ZN(n4638) );
  OAI22_X1 U2248 ( .A1(n4181), .A2(n6299), .B1(n5883), .B2(n6307), .ZN(n4645)
         );
  AOI221_X1 U2249 ( .B1(n6315), .B2(\registers[25][21] ), .C1(n6323), .C2(
        \registers[24][21] ), .A(n4644), .ZN(n4639) );
  OAI22_X1 U2250 ( .A1(n4269), .A2(n6329), .B1(n5965), .B2(n6334), .ZN(n4644)
         );
  AOI221_X1 U2251 ( .B1(\registers[31][22] ), .B2(n6392), .C1(n6394), .C2(
        \registers[30][22] ), .A(n4617), .ZN(n4610) );
  OAI22_X1 U2252 ( .A1(n4201), .A2(n6399), .B1(n5900), .B2(n6409), .ZN(n4617)
         );
  AOI221_X1 U2253 ( .B1(n6282), .B2(\registers[23][22] ), .C1(n6290), .C2(
        \registers[22][22] ), .A(n4625), .ZN(n4618) );
  OAI22_X1 U2254 ( .A1(n4185), .A2(n6298), .B1(n5884), .B2(n6306), .ZN(n4625)
         );
  AOI221_X1 U2255 ( .B1(n6309), .B2(\registers[25][22] ), .C1(n6318), .C2(
        \registers[24][22] ), .A(n4624), .ZN(n4619) );
  OAI22_X1 U2256 ( .A1(n4270), .A2(n6330), .B1(n5966), .B2(n6335), .ZN(n4624)
         );
  AOI221_X1 U2257 ( .B1(\registers[31][23] ), .B2(n4417), .C1(n4418), .C2(
        \registers[30][23] ), .A(n4597), .ZN(n4590) );
  OAI22_X1 U2258 ( .A1(n4203), .A2(n6402), .B1(n5902), .B2(n6405), .ZN(n4597)
         );
  AOI221_X1 U2259 ( .B1(n6283), .B2(\registers[23][23] ), .C1(n6290), .C2(
        \registers[22][23] ), .A(n4605), .ZN(n4598) );
  OAI22_X1 U2260 ( .A1(n4186), .A2(n6299), .B1(n5885), .B2(n6306), .ZN(n4605)
         );
  AOI221_X1 U2261 ( .B1(n6310), .B2(\registers[25][23] ), .C1(n6317), .C2(
        \registers[24][23] ), .A(n4604), .ZN(n4599) );
  OAI22_X1 U2262 ( .A1(n4271), .A2(n6328), .B1(n5967), .B2(n6336), .ZN(n4604)
         );
  AOI221_X1 U2263 ( .B1(\registers[31][24] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][24] ), .A(n4577), .ZN(n4570) );
  OAI22_X1 U2264 ( .A1(n4205), .A2(n6402), .B1(n5904), .B2(n6409), .ZN(n4577)
         );
  AOI221_X1 U2265 ( .B1(n6283), .B2(\registers[23][24] ), .C1(n6291), .C2(
        \registers[22][24] ), .A(n4585), .ZN(n4578) );
  OAI22_X1 U2266 ( .A1(n4187), .A2(n6293), .B1(n5886), .B2(n6304), .ZN(n4585)
         );
  AOI221_X1 U2267 ( .B1(n6310), .B2(\registers[25][24] ), .C1(n6317), .C2(
        \registers[24][24] ), .A(n4584), .ZN(n4579) );
  OAI22_X1 U2268 ( .A1(n4272), .A2(n6331), .B1(n5968), .B2(n6335), .ZN(n4584)
         );
  AOI221_X1 U2269 ( .B1(\registers[31][25] ), .B2(n6392), .C1(n6394), .C2(
        \registers[30][25] ), .A(n4557), .ZN(n4550) );
  OAI22_X1 U2270 ( .A1(n4207), .A2(n6401), .B1(n5906), .B2(n6405), .ZN(n4557)
         );
  AOI221_X1 U2271 ( .B1(n6284), .B2(\registers[23][25] ), .C1(n6289), .C2(
        \registers[22][25] ), .A(n4565), .ZN(n4558) );
  OAI22_X1 U2272 ( .A1(n4188), .A2(n6299), .B1(n5887), .B2(n6307), .ZN(n4565)
         );
  AOI221_X1 U2273 ( .B1(n6311), .B2(\registers[25][25] ), .C1(n6318), .C2(
        \registers[24][25] ), .A(n4564), .ZN(n4559) );
  OAI22_X1 U2274 ( .A1(n4273), .A2(n6325), .B1(n5969), .B2(n6336), .ZN(n4564)
         );
  AOI221_X1 U2275 ( .B1(\registers[31][26] ), .B2(n4417), .C1(n4418), .C2(
        \registers[30][26] ), .A(n4537), .ZN(n4530) );
  OAI22_X1 U2276 ( .A1(n4209), .A2(n6402), .B1(n5908), .B2(n6407), .ZN(n4537)
         );
  AOI221_X1 U2277 ( .B1(n6284), .B2(\registers[23][26] ), .C1(n6291), .C2(
        \registers[22][26] ), .A(n4545), .ZN(n4538) );
  OAI22_X1 U2278 ( .A1(n4189), .A2(n6297), .B1(n5888), .B2(n6302), .ZN(n4545)
         );
  AOI221_X1 U2279 ( .B1(n6311), .B2(\registers[25][26] ), .C1(n6318), .C2(
        \registers[24][26] ), .A(n4544), .ZN(n4539) );
  OAI22_X1 U2280 ( .A1(n4274), .A2(n6331), .B1(n5970), .B2(n6337), .ZN(n4544)
         );
  AOI221_X1 U2281 ( .B1(\registers[31][27] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][27] ), .A(n4517), .ZN(n4510) );
  OAI22_X1 U2282 ( .A1(n4211), .A2(n6399), .B1(n5910), .B2(n6407), .ZN(n4517)
         );
  AOI221_X1 U2283 ( .B1(n6282), .B2(\registers[23][27] ), .C1(n6290), .C2(
        \registers[22][27] ), .A(n4525), .ZN(n4518) );
  OAI22_X1 U2284 ( .A1(n4190), .A2(n6299), .B1(n5889), .B2(n6301), .ZN(n4525)
         );
  AOI221_X1 U2285 ( .B1(n6309), .B2(\registers[25][27] ), .C1(n6321), .C2(
        \registers[24][27] ), .A(n4524), .ZN(n4519) );
  OAI22_X1 U2286 ( .A1(n4275), .A2(n6330), .B1(n5971), .B2(n6338), .ZN(n4524)
         );
  AOI221_X1 U2287 ( .B1(\registers[31][28] ), .B2(n6392), .C1(n6394), .C2(
        \registers[30][28] ), .A(n4497), .ZN(n4490) );
  OAI22_X1 U2288 ( .A1(n4191), .A2(n6398), .B1(n5890), .B2(n6410), .ZN(n4497)
         );
  AOI221_X1 U2289 ( .B1(n6285), .B2(\registers[23][28] ), .C1(n6291), .C2(
        \registers[22][28] ), .A(n4505), .ZN(n4498) );
  OAI22_X1 U2290 ( .A1(n4192), .A2(n6295), .B1(n5891), .B2(n6301), .ZN(n4505)
         );
  AOI221_X1 U2291 ( .B1(n6312), .B2(\registers[25][28] ), .C1(n6317), .C2(
        \registers[24][28] ), .A(n4504), .ZN(n4499) );
  OAI22_X1 U2292 ( .A1(n4276), .A2(n6325), .B1(n5972), .B2(n6333), .ZN(n4504)
         );
  AOI221_X1 U2293 ( .B1(\registers[31][29] ), .B2(n4417), .C1(n4418), .C2(
        \registers[30][29] ), .A(n4477), .ZN(n4470) );
  OAI22_X1 U2294 ( .A1(n4193), .A2(n6397), .B1(n5892), .B2(n6409), .ZN(n4477)
         );
  AOI221_X1 U2295 ( .B1(n6283), .B2(\registers[23][29] ), .C1(n6289), .C2(
        \registers[22][29] ), .A(n4485), .ZN(n4478) );
  OAI22_X1 U2296 ( .A1(n4194), .A2(n6293), .B1(n5893), .B2(n6305), .ZN(n4485)
         );
  AOI221_X1 U2297 ( .B1(n6310), .B2(\registers[25][29] ), .C1(n6319), .C2(
        \registers[24][29] ), .A(n4484), .ZN(n4479) );
  OAI22_X1 U2298 ( .A1(n4277), .A2(n6326), .B1(n5973), .B2(n6334), .ZN(n4484)
         );
  AOI221_X1 U2299 ( .B1(\registers[31][30] ), .B2(n6391), .C1(n6393), .C2(
        \registers[30][30] ), .A(n4457), .ZN(n4450) );
  OAI22_X1 U2300 ( .A1(n4195), .A2(n6400), .B1(n5894), .B2(n6405), .ZN(n4457)
         );
  AOI221_X1 U2301 ( .B1(n6283), .B2(\registers[23][30] ), .C1(n6289), .C2(
        \registers[22][30] ), .A(n4465), .ZN(n4458) );
  OAI22_X1 U2302 ( .A1(n4196), .A2(n6293), .B1(n5895), .B2(n6306), .ZN(n4465)
         );
  AOI221_X1 U2303 ( .B1(n6310), .B2(\registers[25][30] ), .C1(n6319), .C2(
        \registers[24][30] ), .A(n4464), .ZN(n4459) );
  OAI22_X1 U2304 ( .A1(n4278), .A2(n6331), .B1(n5974), .B2(n6337), .ZN(n4464)
         );
  AOI221_X1 U2305 ( .B1(n6392), .B2(\registers[31][31] ), .C1(n6394), .C2(
        \registers[30][31] ), .A(n4419), .ZN(n4398) );
  OAI22_X1 U2306 ( .A1(n4197), .A2(n6401), .B1(n5896), .B2(n6410), .ZN(n4419)
         );
  AOI221_X1 U2307 ( .B1(n6285), .B2(\registers[23][31] ), .C1(n6290), .C2(
        \registers[22][31] ), .A(n4443), .ZN(n4422) );
  OAI22_X1 U2308 ( .A1(n4198), .A2(n6298), .B1(n5897), .B2(n6306), .ZN(n4443)
         );
  AOI221_X1 U2309 ( .B1(n6312), .B2(\registers[25][31] ), .C1(n6320), .C2(
        \registers[24][31] ), .A(n4438), .ZN(n4423) );
  OAI22_X1 U2310 ( .A1(n4279), .A2(n6325), .B1(n5975), .B2(n6338), .ZN(n4438)
         );
  NOR3_X1 U2311 ( .A1(n5757), .A2(n2720), .A3(n5758), .ZN(n5756) );
  XNOR2_X1 U2312 ( .A(n1857), .B(add_rd1[2]), .ZN(n5757) );
  XNOR2_X1 U2313 ( .A(add_wr[4]), .B(n5748), .ZN(n5758) );
  NOR3_X1 U2314 ( .A1(n5089), .A2(n2720), .A3(n5090), .ZN(n5088) );
  XNOR2_X1 U2315 ( .A(n1857), .B(add_rd2[2]), .ZN(n5089) );
  XNOR2_X1 U2316 ( .A(add_wr[4]), .B(n5081), .ZN(n5090) );
  AND3_X1 U2317 ( .A1(n1859), .A2(n1858), .A3(add_wr[2]), .ZN(n1894) );
  OR3_X1 U2318 ( .A1(rd1), .A2(n5752), .A3(n2719), .ZN(n6073) );
  OR3_X1 U2319 ( .A1(rd1), .A2(n5752), .A3(n2719), .ZN(n5091) );
  OR3_X1 U2320 ( .A1(rd2), .A2(n5084), .A3(n2719), .ZN(n6278) );
  OR3_X1 U2321 ( .A1(rd2), .A2(n5084), .A3(n2719), .ZN(n4392) );
  OR3_X1 U2322 ( .A1(rd1), .A2(n5752), .A3(n2719), .ZN(n6072) );
  OR3_X1 U2323 ( .A1(rd2), .A2(n5084), .A3(n2719), .ZN(n6277) );
  INV_X1 U2324 ( .A(add_rd1[4]), .ZN(n5748) );
  INV_X1 U2325 ( .A(add_wr[2]), .ZN(n1857) );
  INV_X1 U2326 ( .A(add_rd1[0]), .ZN(n5745) );
  INV_X1 U2327 ( .A(add_rd1[3]), .ZN(n5744) );
  AND3_X1 U2328 ( .A1(add_wr[3]), .A2(add_wr[2]), .A3(n2858), .ZN(n4319) );
  AND3_X1 U2329 ( .A1(add_wr[3]), .A2(n1857), .A3(n2858), .ZN(n4182) );
  AND3_X1 U2330 ( .A1(add_wr[2]), .A2(n1859), .A3(add_wr[3]), .ZN(n2616) );
  AND3_X1 U2331 ( .A1(n1859), .A2(n1857), .A3(add_wr[3]), .ZN(n2031) );
  AND3_X1 U2332 ( .A1(add_wr[2]), .A2(n1858), .A3(n2858), .ZN(n2893) );
  NAND4_X1 U2333 ( .A1(n5753), .A2(n5754), .A3(n5755), .A4(n5756), .ZN(n5718)
         );
  XNOR2_X1 U2334 ( .A(add_rd1[3]), .B(add_wr[3]), .ZN(n5753) );
  XNOR2_X1 U2335 ( .A(add_rd1[1]), .B(add_wr[1]), .ZN(n5754) );
  XNOR2_X1 U2336 ( .A(add_wr[0]), .B(add_rd1[0]), .ZN(n5755) );
  NAND4_X1 U2337 ( .A1(n5085), .A2(n5086), .A3(n5087), .A4(n5088), .ZN(n5050)
         );
  XNOR2_X1 U2338 ( .A(add_rd2[1]), .B(add_wr[1]), .ZN(n5086) );
  XNOR2_X1 U2339 ( .A(add_rd2[3]), .B(add_wr[3]), .ZN(n5085) );
  XNOR2_X1 U2340 ( .A(add_wr[0]), .B(add_rd2[0]), .ZN(n5087) );
  AND3_X1 U2341 ( .A1(n6072), .A2(n5718), .A3(enable), .ZN(n5096) );
  AND3_X1 U2342 ( .A1(n6277), .A2(n5050), .A3(enable), .ZN(n4397) );
  AND3_X1 U2343 ( .A1(wr), .A2(enable), .A3(add_wr[4]), .ZN(n2858) );
  INV_X1 U2344 ( .A(wr), .ZN(n2720) );
  INV_X1 U2345 ( .A(add_wr[3]), .ZN(n1858) );
  INV_X1 U2346 ( .A(add_rd1[2]), .ZN(n5749) );
  INV_X1 U2347 ( .A(add_rd1[1]), .ZN(n5751) );
  INV_X1 U2348 ( .A(add_wr[0]), .ZN(n4354) );
  AOI221_X1 U2349 ( .B1(n5116), .B2(\registers[31][20] ), .C1(n5117), .C2(
        \registers[30][20] ), .A(n5345), .ZN(n5338) );
  OAI22_X1 U2350 ( .A1(n4199), .A2(n6187), .B1(n5898), .B2(n6199), .ZN(n5345)
         );
  AOI221_X1 U2351 ( .B1(n6182), .B2(\registers[31][21] ), .C1(n6184), .C2(
        \registers[30][21] ), .A(n5326), .ZN(n5319) );
  OAI22_X1 U2352 ( .A1(n4200), .A2(n6188), .B1(n5899), .B2(n6201), .ZN(n5326)
         );
  AOI221_X1 U2353 ( .B1(n6183), .B2(\registers[31][22] ), .C1(n6185), .C2(
        \registers[30][22] ), .A(n5307), .ZN(n5300) );
  OAI22_X1 U2354 ( .A1(n4201), .A2(n6192), .B1(n5900), .B2(n6200), .ZN(n5307)
         );
  AOI221_X1 U2355 ( .B1(n6136), .B2(\registers[6][22] ), .C1(n6144), .C2(
        \registers[7][22] ), .A(n5313), .ZN(n5310) );
  OAI22_X1 U2356 ( .A1(n4202), .A2(n6147), .B1(n5901), .B2(n6160), .ZN(n5313)
         );
  AOI221_X1 U2357 ( .B1(n5116), .B2(\registers[31][23] ), .C1(n5117), .C2(
        \registers[30][23] ), .A(n5288), .ZN(n5281) );
  OAI22_X1 U2358 ( .A1(n4203), .A2(n6188), .B1(n5902), .B2(n6201), .ZN(n5288)
         );
  AOI221_X1 U2359 ( .B1(n6138), .B2(\registers[6][23] ), .C1(n6144), .C2(
        \registers[7][23] ), .A(n5294), .ZN(n5291) );
  OAI22_X1 U2360 ( .A1(n4204), .A2(n6153), .B1(n5903), .B2(n6155), .ZN(n5294)
         );
  AOI221_X1 U2361 ( .B1(n6182), .B2(\registers[31][24] ), .C1(n6184), .C2(
        \registers[30][24] ), .A(n5269), .ZN(n5262) );
  OAI22_X1 U2362 ( .A1(n4205), .A2(n6193), .B1(n5904), .B2(n6201), .ZN(n5269)
         );
  AOI221_X1 U2363 ( .B1(n6139), .B2(\registers[6][24] ), .C1(n6145), .C2(
        \registers[7][24] ), .A(n5275), .ZN(n5272) );
  OAI22_X1 U2364 ( .A1(n4206), .A2(n6147), .B1(n5905), .B2(n6161), .ZN(n5275)
         );
  AOI221_X1 U2365 ( .B1(n6183), .B2(\registers[31][25] ), .C1(n6185), .C2(
        \registers[30][25] ), .A(n5250), .ZN(n5243) );
  OAI22_X1 U2366 ( .A1(n4207), .A2(n6192), .B1(n5906), .B2(n6195), .ZN(n5250)
         );
  AOI221_X1 U2367 ( .B1(n6137), .B2(\registers[6][25] ), .C1(n6143), .C2(
        \registers[7][25] ), .A(n5256), .ZN(n5253) );
  OAI22_X1 U2368 ( .A1(n4208), .A2(n6152), .B1(n5907), .B2(n6159), .ZN(n5256)
         );
  AOI221_X1 U2369 ( .B1(n5116), .B2(\registers[31][26] ), .C1(n5117), .C2(
        \registers[30][26] ), .A(n5231), .ZN(n5224) );
  OAI22_X1 U2370 ( .A1(n4209), .A2(n6193), .B1(n5908), .B2(n6200), .ZN(n5231)
         );
  AOI221_X1 U2371 ( .B1(n6140), .B2(\registers[6][26] ), .C1(n6145), .C2(
        \registers[7][26] ), .A(n5237), .ZN(n5234) );
  OAI22_X1 U2372 ( .A1(n4210), .A2(n6152), .B1(n5909), .B2(n6161), .ZN(n5237)
         );
  AOI221_X1 U2373 ( .B1(n6182), .B2(\registers[31][27] ), .C1(n6184), .C2(
        \registers[30][27] ), .A(n5212), .ZN(n5205) );
  OAI22_X1 U2374 ( .A1(n4211), .A2(n6187), .B1(n5910), .B2(n6199), .ZN(n5212)
         );
  AOI221_X1 U2375 ( .B1(n6140), .B2(\registers[6][27] ), .C1(n6144), .C2(
        \registers[7][27] ), .A(n5218), .ZN(n5215) );
  OAI22_X1 U2376 ( .A1(n4212), .A2(n6147), .B1(n5911), .B2(n6155), .ZN(n5218)
         );
  AOI221_X1 U2377 ( .B1(n6203), .B2(\registers[21][22] ), .C1(n6215), .C2(
        \registers[20][22] ), .A(n5306), .ZN(n5301) );
  OAI22_X1 U2378 ( .A1(n4213), .A2(n6219), .B1(n5912), .B2(n6227), .ZN(n5306)
         );
  AOI221_X1 U2379 ( .B1(n6109), .B2(\registers[29][22] ), .C1(n6117), .C2(
        \registers[28][22] ), .A(n5314), .ZN(n5309) );
  OAI22_X1 U2380 ( .A1(n4280), .A2(n6125), .B1(n5976), .B2(n6128), .ZN(n5314)
         );
  AOI221_X1 U2381 ( .B1(n6204), .B2(\registers[21][23] ), .C1(n6211), .C2(
        \registers[20][23] ), .A(n5287), .ZN(n5282) );
  OAI22_X1 U2382 ( .A1(n4214), .A2(n6225), .B1(n5913), .B2(n6233), .ZN(n5287)
         );
  AOI221_X1 U2383 ( .B1(n6111), .B2(\registers[29][23] ), .C1(n6117), .C2(
        \registers[28][23] ), .A(n5295), .ZN(n5290) );
  OAI22_X1 U2384 ( .A1(n4281), .A2(n6124), .B1(n5977), .B2(n6132), .ZN(n5295)
         );
  AOI221_X1 U2385 ( .B1(n6203), .B2(\registers[21][24] ), .C1(n6214), .C2(
        \registers[20][24] ), .A(n5268), .ZN(n5263) );
  OAI22_X1 U2386 ( .A1(n4215), .A2(n6219), .B1(n5914), .B2(n6233), .ZN(n5268)
         );
  AOI221_X1 U2387 ( .B1(n6112), .B2(\registers[29][24] ), .C1(n6118), .C2(
        \registers[28][24] ), .A(n5276), .ZN(n5271) );
  OAI22_X1 U2388 ( .A1(n4282), .A2(n6120), .B1(n5978), .B2(n6134), .ZN(n5276)
         );
  AOI221_X1 U2389 ( .B1(n6205), .B2(\registers[21][25] ), .C1(n6212), .C2(
        \registers[20][25] ), .A(n5249), .ZN(n5244) );
  OAI22_X1 U2390 ( .A1(n4216), .A2(n6224), .B1(n5915), .B2(n6232), .ZN(n5249)
         );
  AOI221_X1 U2391 ( .B1(n6110), .B2(\registers[29][25] ), .C1(n6116), .C2(
        \registers[28][25] ), .A(n5257), .ZN(n5252) );
  OAI22_X1 U2392 ( .A1(n4283), .A2(n6120), .B1(n5979), .B2(n6133), .ZN(n5257)
         );
  AOI221_X1 U2393 ( .B1(n6204), .B2(\registers[21][26] ), .C1(n6217), .C2(
        \registers[20][26] ), .A(n5230), .ZN(n5225) );
  OAI22_X1 U2394 ( .A1(n4218), .A2(n6220), .B1(n5916), .B2(n6232), .ZN(n5230)
         );
  AOI221_X1 U2395 ( .B1(n6113), .B2(\registers[29][26] ), .C1(n6118), .C2(
        \registers[28][26] ), .A(n5238), .ZN(n5233) );
  OAI22_X1 U2396 ( .A1(n4284), .A2(n6124), .B1(n5980), .B2(n6131), .ZN(n5238)
         );
  AOI221_X1 U2397 ( .B1(n6207), .B2(\registers[21][27] ), .C1(n6212), .C2(
        \registers[20][27] ), .A(n5211), .ZN(n5206) );
  OAI22_X1 U2398 ( .A1(n4219), .A2(n6225), .B1(n5917), .B2(n6228), .ZN(n5211)
         );
  AOI221_X1 U2399 ( .B1(n6113), .B2(\registers[29][27] ), .C1(n6117), .C2(
        \registers[28][27] ), .A(n5219), .ZN(n5214) );
  OAI22_X1 U2400 ( .A1(n4287), .A2(n6126), .B1(n5981), .B2(n6132), .ZN(n5219)
         );
  INV_X1 U2401 ( .A(n5046), .ZN(n3084) );
  AOI22_X1 U2402 ( .A1(datain[0]), .A2(n5982), .B1(n6493), .B2(
        \registers[31][0] ), .ZN(n5046) );
  INV_X1 U2403 ( .A(n5026), .ZN(n3086) );
  AOI22_X1 U2404 ( .A1(datain[1]), .A2(n5982), .B1(n6494), .B2(
        \registers[31][1] ), .ZN(n5026) );
  INV_X1 U2405 ( .A(n5006), .ZN(n3088) );
  AOI22_X1 U2406 ( .A1(datain[2]), .A2(n5982), .B1(n6495), .B2(
        \registers[31][2] ), .ZN(n5006) );
  INV_X1 U2407 ( .A(n4986), .ZN(n3090) );
  AOI22_X1 U2408 ( .A1(datain[3]), .A2(n5982), .B1(n6498), .B2(
        \registers[31][3] ), .ZN(n4986) );
  INV_X1 U2409 ( .A(n4966), .ZN(n3092) );
  AOI22_X1 U2410 ( .A1(datain[4]), .A2(n5982), .B1(n6494), .B2(
        \registers[31][4] ), .ZN(n4966) );
  INV_X1 U2411 ( .A(n4946), .ZN(n3094) );
  AOI22_X1 U2412 ( .A1(datain[5]), .A2(n5982), .B1(n6495), .B2(
        \registers[31][5] ), .ZN(n4946) );
  INV_X1 U2413 ( .A(n4926), .ZN(n3096) );
  AOI22_X1 U2414 ( .A1(datain[6]), .A2(n5982), .B1(n6495), .B2(
        \registers[31][6] ), .ZN(n4926) );
  INV_X1 U2415 ( .A(n4906), .ZN(n3098) );
  AOI22_X1 U2416 ( .A1(datain[7]), .A2(n5982), .B1(n6496), .B2(
        \registers[31][7] ), .ZN(n4906) );
  INV_X1 U2417 ( .A(n4886), .ZN(n3100) );
  AOI22_X1 U2418 ( .A1(datain[8]), .A2(n5982), .B1(n6496), .B2(
        \registers[31][8] ), .ZN(n4886) );
  INV_X1 U2419 ( .A(n4866), .ZN(n3102) );
  AOI22_X1 U2420 ( .A1(datain[9]), .A2(n5982), .B1(n6497), .B2(
        \registers[31][9] ), .ZN(n4866) );
  INV_X1 U2421 ( .A(n4846), .ZN(n3104) );
  AOI22_X1 U2422 ( .A1(datain[10]), .A2(n5982), .B1(n6497), .B2(
        \registers[31][10] ), .ZN(n4846) );
  INV_X1 U2423 ( .A(n4826), .ZN(n3106) );
  AOI22_X1 U2424 ( .A1(datain[11]), .A2(n5982), .B1(n6499), .B2(
        \registers[31][11] ), .ZN(n4826) );
  INV_X1 U2425 ( .A(n4806), .ZN(n3108) );
  AOI22_X1 U2426 ( .A1(datain[12]), .A2(n5983), .B1(n6493), .B2(
        \registers[31][12] ), .ZN(n4806) );
  INV_X1 U2427 ( .A(n4786), .ZN(n3110) );
  AOI22_X1 U2428 ( .A1(datain[13]), .A2(n5983), .B1(n6494), .B2(
        \registers[31][13] ), .ZN(n4786) );
  INV_X1 U2429 ( .A(n4766), .ZN(n3112) );
  AOI22_X1 U2430 ( .A1(datain[14]), .A2(n5983), .B1(n6495), .B2(
        \registers[31][14] ), .ZN(n4766) );
  INV_X1 U2431 ( .A(n4746), .ZN(n3114) );
  AOI22_X1 U2432 ( .A1(datain[15]), .A2(n5983), .B1(n6494), .B2(
        \registers[31][15] ), .ZN(n4746) );
  INV_X1 U2433 ( .A(n4726), .ZN(n3116) );
  AOI22_X1 U2434 ( .A1(datain[16]), .A2(n5983), .B1(n6496), .B2(
        \registers[31][16] ), .ZN(n4726) );
  INV_X1 U2435 ( .A(n4706), .ZN(n3118) );
  AOI22_X1 U2436 ( .A1(datain[17]), .A2(n5983), .B1(n6496), .B2(
        \registers[31][17] ), .ZN(n4706) );
  INV_X1 U2437 ( .A(n4686), .ZN(n3120) );
  AOI22_X1 U2438 ( .A1(datain[18]), .A2(n5983), .B1(n6497), .B2(
        \registers[31][18] ), .ZN(n4686) );
  INV_X1 U2439 ( .A(n4666), .ZN(n3122) );
  AOI22_X1 U2440 ( .A1(datain[19]), .A2(n5983), .B1(n6496), .B2(
        \registers[31][19] ), .ZN(n4666) );
  INV_X1 U2441 ( .A(n4646), .ZN(n3124) );
  AOI22_X1 U2442 ( .A1(datain[20]), .A2(n5983), .B1(n6498), .B2(
        \registers[31][20] ), .ZN(n4646) );
  INV_X1 U2443 ( .A(n4626), .ZN(n3126) );
  AOI22_X1 U2444 ( .A1(datain[21]), .A2(n5983), .B1(n6499), .B2(
        \registers[31][21] ), .ZN(n4626) );
  INV_X1 U2445 ( .A(n4606), .ZN(n3128) );
  AOI22_X1 U2446 ( .A1(datain[22]), .A2(n5983), .B1(n6498), .B2(
        \registers[31][22] ), .ZN(n4606) );
  INV_X1 U2447 ( .A(n4586), .ZN(n3130) );
  AOI22_X1 U2448 ( .A1(datain[23]), .A2(n5983), .B1(n6498), .B2(
        \registers[31][23] ), .ZN(n4586) );
  INV_X1 U2449 ( .A(n4566), .ZN(n3132) );
  AOI22_X1 U2450 ( .A1(datain[24]), .A2(n5984), .B1(n6499), .B2(
        \registers[31][24] ), .ZN(n4566) );
  INV_X1 U2451 ( .A(n4546), .ZN(n3134) );
  AOI22_X1 U2452 ( .A1(datain[25]), .A2(n5984), .B1(n6499), .B2(
        \registers[31][25] ), .ZN(n4546) );
  INV_X1 U2453 ( .A(n4526), .ZN(n3136) );
  AOI22_X1 U2454 ( .A1(datain[26]), .A2(n5984), .B1(n6493), .B2(
        \registers[31][26] ), .ZN(n4526) );
  INV_X1 U2455 ( .A(n4506), .ZN(n3138) );
  AOI22_X1 U2456 ( .A1(datain[27]), .A2(n5984), .B1(n6493), .B2(
        \registers[31][27] ), .ZN(n4506) );
  INV_X1 U2457 ( .A(n4486), .ZN(n3140) );
  AOI22_X1 U2458 ( .A1(datain[28]), .A2(n5984), .B1(n6493), .B2(
        \registers[31][28] ), .ZN(n4486) );
  INV_X1 U2459 ( .A(n4466), .ZN(n3142) );
  AOI22_X1 U2460 ( .A1(datain[29]), .A2(n5984), .B1(n6499), .B2(
        \registers[31][29] ), .ZN(n4466) );
  INV_X1 U2461 ( .A(n4446), .ZN(n3144) );
  AOI22_X1 U2462 ( .A1(datain[30]), .A2(n5984), .B1(n6494), .B2(
        \registers[31][30] ), .ZN(n4446) );
  INV_X1 U2463 ( .A(n4389), .ZN(n3146) );
  AOI22_X1 U2464 ( .A1(datain[31]), .A2(n5984), .B1(n6497), .B2(
        \registers[31][31] ), .ZN(n4389) );
  INV_X1 U2465 ( .A(n4388), .ZN(n3147) );
  AOI22_X1 U2466 ( .A1(datain[0]), .A2(n5985), .B1(n6502), .B2(
        \registers[30][0] ), .ZN(n4388) );
  INV_X1 U2467 ( .A(n4387), .ZN(n3148) );
  AOI22_X1 U2468 ( .A1(datain[1]), .A2(n5985), .B1(n6503), .B2(
        \registers[30][1] ), .ZN(n4387) );
  INV_X1 U2469 ( .A(n4386), .ZN(n3149) );
  AOI22_X1 U2470 ( .A1(datain[2]), .A2(n5985), .B1(n6504), .B2(
        \registers[30][2] ), .ZN(n4386) );
  INV_X1 U2471 ( .A(n4385), .ZN(n3150) );
  AOI22_X1 U2472 ( .A1(datain[3]), .A2(n5985), .B1(n6507), .B2(
        \registers[30][3] ), .ZN(n4385) );
  INV_X1 U2473 ( .A(n4384), .ZN(n3151) );
  AOI22_X1 U2474 ( .A1(datain[4]), .A2(n5985), .B1(n6503), .B2(
        \registers[30][4] ), .ZN(n4384) );
  INV_X1 U2475 ( .A(n4383), .ZN(n3152) );
  AOI22_X1 U2476 ( .A1(datain[5]), .A2(n5985), .B1(n6504), .B2(
        \registers[30][5] ), .ZN(n4383) );
  INV_X1 U2477 ( .A(n4382), .ZN(n3153) );
  AOI22_X1 U2478 ( .A1(datain[6]), .A2(n5985), .B1(n6504), .B2(
        \registers[30][6] ), .ZN(n4382) );
  INV_X1 U2479 ( .A(n4381), .ZN(n3154) );
  AOI22_X1 U2480 ( .A1(datain[7]), .A2(n5985), .B1(n6505), .B2(
        \registers[30][7] ), .ZN(n4381) );
  INV_X1 U2481 ( .A(n4380), .ZN(n3155) );
  AOI22_X1 U2482 ( .A1(datain[8]), .A2(n5985), .B1(n6505), .B2(
        \registers[30][8] ), .ZN(n4380) );
  INV_X1 U2483 ( .A(n4379), .ZN(n3156) );
  AOI22_X1 U2484 ( .A1(datain[9]), .A2(n5985), .B1(n6506), .B2(
        \registers[30][9] ), .ZN(n4379) );
  INV_X1 U2485 ( .A(n4378), .ZN(n3157) );
  AOI22_X1 U2486 ( .A1(datain[10]), .A2(n5985), .B1(n6506), .B2(
        \registers[30][10] ), .ZN(n4378) );
  INV_X1 U2487 ( .A(n4377), .ZN(n3158) );
  AOI22_X1 U2488 ( .A1(datain[11]), .A2(n5985), .B1(n6508), .B2(
        \registers[30][11] ), .ZN(n4377) );
  INV_X1 U2489 ( .A(n4376), .ZN(n3159) );
  AOI22_X1 U2490 ( .A1(datain[12]), .A2(n5986), .B1(n6502), .B2(
        \registers[30][12] ), .ZN(n4376) );
  INV_X1 U2491 ( .A(n4375), .ZN(n3160) );
  AOI22_X1 U2492 ( .A1(datain[13]), .A2(n5986), .B1(n6503), .B2(
        \registers[30][13] ), .ZN(n4375) );
  INV_X1 U2493 ( .A(n4374), .ZN(n3161) );
  AOI22_X1 U2494 ( .A1(datain[14]), .A2(n5986), .B1(n6504), .B2(
        \registers[30][14] ), .ZN(n4374) );
  INV_X1 U2495 ( .A(n4373), .ZN(n3162) );
  AOI22_X1 U2496 ( .A1(datain[15]), .A2(n5986), .B1(n6503), .B2(
        \registers[30][15] ), .ZN(n4373) );
  INV_X1 U2497 ( .A(n4372), .ZN(n3163) );
  AOI22_X1 U2498 ( .A1(datain[16]), .A2(n5986), .B1(n6505), .B2(
        \registers[30][16] ), .ZN(n4372) );
  INV_X1 U2499 ( .A(n4371), .ZN(n3164) );
  AOI22_X1 U2500 ( .A1(datain[17]), .A2(n5986), .B1(n6505), .B2(
        \registers[30][17] ), .ZN(n4371) );
  INV_X1 U2501 ( .A(n4370), .ZN(n3165) );
  AOI22_X1 U2502 ( .A1(datain[18]), .A2(n5986), .B1(n6506), .B2(
        \registers[30][18] ), .ZN(n4370) );
  INV_X1 U2503 ( .A(n4369), .ZN(n3166) );
  AOI22_X1 U2504 ( .A1(datain[19]), .A2(n5986), .B1(n6505), .B2(
        \registers[30][19] ), .ZN(n4369) );
  INV_X1 U2505 ( .A(n4368), .ZN(n3167) );
  AOI22_X1 U2506 ( .A1(datain[20]), .A2(n5986), .B1(n6507), .B2(
        \registers[30][20] ), .ZN(n4368) );
  INV_X1 U2507 ( .A(n4367), .ZN(n3168) );
  AOI22_X1 U2508 ( .A1(datain[21]), .A2(n5986), .B1(n6508), .B2(
        \registers[30][21] ), .ZN(n4367) );
  INV_X1 U2509 ( .A(n4366), .ZN(n3169) );
  AOI22_X1 U2510 ( .A1(datain[22]), .A2(n5986), .B1(n6507), .B2(
        \registers[30][22] ), .ZN(n4366) );
  INV_X1 U2511 ( .A(n4365), .ZN(n3170) );
  AOI22_X1 U2512 ( .A1(datain[23]), .A2(n5986), .B1(n6507), .B2(
        \registers[30][23] ), .ZN(n4365) );
  INV_X1 U2513 ( .A(n4364), .ZN(n3171) );
  AOI22_X1 U2514 ( .A1(datain[24]), .A2(n5987), .B1(n6508), .B2(
        \registers[30][24] ), .ZN(n4364) );
  INV_X1 U2515 ( .A(n4363), .ZN(n3172) );
  AOI22_X1 U2516 ( .A1(datain[25]), .A2(n5987), .B1(n6508), .B2(
        \registers[30][25] ), .ZN(n4363) );
  INV_X1 U2517 ( .A(n4362), .ZN(n3173) );
  AOI22_X1 U2518 ( .A1(datain[26]), .A2(n5987), .B1(n6502), .B2(
        \registers[30][26] ), .ZN(n4362) );
  INV_X1 U2519 ( .A(n4361), .ZN(n3174) );
  AOI22_X1 U2520 ( .A1(datain[27]), .A2(n5987), .B1(n6502), .B2(
        \registers[30][27] ), .ZN(n4361) );
  INV_X1 U2521 ( .A(n4360), .ZN(n3175) );
  AOI22_X1 U2522 ( .A1(datain[28]), .A2(n5987), .B1(n6502), .B2(
        \registers[30][28] ), .ZN(n4360) );
  INV_X1 U2523 ( .A(n4359), .ZN(n3176) );
  AOI22_X1 U2524 ( .A1(datain[29]), .A2(n5987), .B1(n6508), .B2(
        \registers[30][29] ), .ZN(n4359) );
  INV_X1 U2525 ( .A(n4358), .ZN(n3177) );
  AOI22_X1 U2526 ( .A1(datain[30]), .A2(n5987), .B1(n6503), .B2(
        \registers[30][30] ), .ZN(n4358) );
  INV_X1 U2527 ( .A(n4355), .ZN(n3178) );
  AOI22_X1 U2528 ( .A1(datain[31]), .A2(n5987), .B1(n6506), .B2(
        \registers[30][31] ), .ZN(n4355) );
  INV_X1 U2529 ( .A(n4147), .ZN(n3371) );
  AOI22_X1 U2530 ( .A1(datain[0]), .A2(n6006), .B1(n6560), .B2(
        \registers[23][0] ), .ZN(n4147) );
  INV_X1 U2531 ( .A(n4146), .ZN(n3372) );
  AOI22_X1 U2532 ( .A1(datain[1]), .A2(n6006), .B1(n6561), .B2(
        \registers[23][1] ), .ZN(n4146) );
  INV_X1 U2533 ( .A(n4145), .ZN(n3373) );
  AOI22_X1 U2534 ( .A1(datain[2]), .A2(n6006), .B1(n6562), .B2(
        \registers[23][2] ), .ZN(n4145) );
  INV_X1 U2535 ( .A(n4144), .ZN(n3374) );
  AOI22_X1 U2536 ( .A1(datain[3]), .A2(n6006), .B1(n6565), .B2(
        \registers[23][3] ), .ZN(n4144) );
  INV_X1 U2537 ( .A(n4143), .ZN(n3375) );
  AOI22_X1 U2538 ( .A1(datain[4]), .A2(n6006), .B1(n6561), .B2(
        \registers[23][4] ), .ZN(n4143) );
  INV_X1 U2539 ( .A(n4142), .ZN(n3376) );
  AOI22_X1 U2540 ( .A1(datain[5]), .A2(n6006), .B1(n6562), .B2(
        \registers[23][5] ), .ZN(n4142) );
  INV_X1 U2541 ( .A(n4141), .ZN(n3377) );
  AOI22_X1 U2542 ( .A1(datain[6]), .A2(n6006), .B1(n6562), .B2(
        \registers[23][6] ), .ZN(n4141) );
  INV_X1 U2543 ( .A(n4140), .ZN(n3378) );
  AOI22_X1 U2544 ( .A1(datain[7]), .A2(n6006), .B1(n6563), .B2(
        \registers[23][7] ), .ZN(n4140) );
  INV_X1 U2545 ( .A(n4139), .ZN(n3379) );
  AOI22_X1 U2546 ( .A1(datain[8]), .A2(n6006), .B1(n6563), .B2(
        \registers[23][8] ), .ZN(n4139) );
  INV_X1 U2547 ( .A(n3017), .ZN(n3380) );
  AOI22_X1 U2548 ( .A1(datain[9]), .A2(n6006), .B1(n6564), .B2(
        \registers[23][9] ), .ZN(n3017) );
  INV_X1 U2549 ( .A(n3015), .ZN(n3381) );
  AOI22_X1 U2550 ( .A1(datain[10]), .A2(n6006), .B1(n6564), .B2(
        \registers[23][10] ), .ZN(n3015) );
  INV_X1 U2551 ( .A(n3013), .ZN(n3382) );
  AOI22_X1 U2552 ( .A1(datain[11]), .A2(n6006), .B1(n6566), .B2(
        \registers[23][11] ), .ZN(n3013) );
  INV_X1 U2553 ( .A(n3011), .ZN(n3383) );
  AOI22_X1 U2554 ( .A1(datain[12]), .A2(n6007), .B1(n6560), .B2(
        \registers[23][12] ), .ZN(n3011) );
  INV_X1 U2555 ( .A(n3009), .ZN(n3384) );
  AOI22_X1 U2556 ( .A1(datain[13]), .A2(n6007), .B1(n6561), .B2(
        \registers[23][13] ), .ZN(n3009) );
  INV_X1 U2557 ( .A(n3007), .ZN(n3385) );
  AOI22_X1 U2558 ( .A1(datain[14]), .A2(n6007), .B1(n6562), .B2(
        \registers[23][14] ), .ZN(n3007) );
  INV_X1 U2559 ( .A(n3005), .ZN(n3386) );
  AOI22_X1 U2560 ( .A1(datain[15]), .A2(n6007), .B1(n6561), .B2(
        \registers[23][15] ), .ZN(n3005) );
  INV_X1 U2561 ( .A(n3003), .ZN(n3387) );
  AOI22_X1 U2562 ( .A1(datain[16]), .A2(n6007), .B1(n6563), .B2(
        \registers[23][16] ), .ZN(n3003) );
  INV_X1 U2563 ( .A(n3001), .ZN(n3388) );
  AOI22_X1 U2564 ( .A1(datain[17]), .A2(n6007), .B1(n6563), .B2(
        \registers[23][17] ), .ZN(n3001) );
  INV_X1 U2565 ( .A(n2999), .ZN(n3389) );
  AOI22_X1 U2566 ( .A1(datain[18]), .A2(n6007), .B1(n6564), .B2(
        \registers[23][18] ), .ZN(n2999) );
  INV_X1 U2567 ( .A(n2997), .ZN(n3390) );
  AOI22_X1 U2568 ( .A1(datain[19]), .A2(n6007), .B1(n6563), .B2(
        \registers[23][19] ), .ZN(n2997) );
  INV_X1 U2569 ( .A(n2995), .ZN(n3391) );
  AOI22_X1 U2570 ( .A1(datain[20]), .A2(n6007), .B1(n6565), .B2(
        \registers[23][20] ), .ZN(n2995) );
  INV_X1 U2571 ( .A(n2993), .ZN(n3392) );
  AOI22_X1 U2572 ( .A1(datain[21]), .A2(n6007), .B1(n6566), .B2(
        \registers[23][21] ), .ZN(n2993) );
  INV_X1 U2573 ( .A(n2991), .ZN(n3393) );
  AOI22_X1 U2574 ( .A1(datain[22]), .A2(n6007), .B1(n6565), .B2(
        \registers[23][22] ), .ZN(n2991) );
  INV_X1 U2575 ( .A(n2989), .ZN(n3394) );
  AOI22_X1 U2576 ( .A1(datain[23]), .A2(n6007), .B1(n6565), .B2(
        \registers[23][23] ), .ZN(n2989) );
  INV_X1 U2577 ( .A(n2987), .ZN(n3395) );
  AOI22_X1 U2578 ( .A1(datain[24]), .A2(n6008), .B1(n6566), .B2(
        \registers[23][24] ), .ZN(n2987) );
  INV_X1 U2579 ( .A(n2985), .ZN(n3396) );
  AOI22_X1 U2580 ( .A1(datain[25]), .A2(n6008), .B1(n6566), .B2(
        \registers[23][25] ), .ZN(n2985) );
  INV_X1 U2581 ( .A(n2983), .ZN(n3397) );
  AOI22_X1 U2582 ( .A1(datain[26]), .A2(n6008), .B1(n6560), .B2(
        \registers[23][26] ), .ZN(n2983) );
  INV_X1 U2583 ( .A(n2981), .ZN(n3398) );
  AOI22_X1 U2584 ( .A1(datain[27]), .A2(n6008), .B1(n6560), .B2(
        \registers[23][27] ), .ZN(n2981) );
  INV_X1 U2585 ( .A(n2979), .ZN(n3399) );
  AOI22_X1 U2586 ( .A1(datain[28]), .A2(n6008), .B1(n6560), .B2(
        \registers[23][28] ), .ZN(n2979) );
  INV_X1 U2587 ( .A(n2977), .ZN(n3400) );
  AOI22_X1 U2588 ( .A1(datain[29]), .A2(n6008), .B1(n6566), .B2(
        \registers[23][29] ), .ZN(n2977) );
  INV_X1 U2589 ( .A(n2975), .ZN(n3401) );
  AOI22_X1 U2590 ( .A1(datain[30]), .A2(n6008), .B1(n6561), .B2(
        \registers[23][30] ), .ZN(n2975) );
  INV_X1 U2591 ( .A(n2969), .ZN(n3402) );
  AOI22_X1 U2592 ( .A1(datain[31]), .A2(n6008), .B1(n6564), .B2(
        \registers[23][31] ), .ZN(n2969) );
  INV_X1 U2593 ( .A(n2967), .ZN(n3403) );
  AOI22_X1 U2594 ( .A1(datain[0]), .A2(n6009), .B1(n6569), .B2(
        \registers[22][0] ), .ZN(n2967) );
  INV_X1 U2595 ( .A(n2965), .ZN(n3404) );
  AOI22_X1 U2596 ( .A1(datain[1]), .A2(n6009), .B1(n6570), .B2(
        \registers[22][1] ), .ZN(n2965) );
  INV_X1 U2597 ( .A(n2963), .ZN(n3405) );
  AOI22_X1 U2598 ( .A1(datain[2]), .A2(n6009), .B1(n6571), .B2(
        \registers[22][2] ), .ZN(n2963) );
  INV_X1 U2599 ( .A(n2961), .ZN(n3406) );
  AOI22_X1 U2600 ( .A1(datain[3]), .A2(n6009), .B1(n6574), .B2(
        \registers[22][3] ), .ZN(n2961) );
  INV_X1 U2601 ( .A(n2959), .ZN(n3407) );
  AOI22_X1 U2602 ( .A1(datain[4]), .A2(n6009), .B1(n6570), .B2(
        \registers[22][4] ), .ZN(n2959) );
  INV_X1 U2603 ( .A(n2957), .ZN(n3408) );
  AOI22_X1 U2604 ( .A1(datain[5]), .A2(n6009), .B1(n6571), .B2(
        \registers[22][5] ), .ZN(n2957) );
  INV_X1 U2605 ( .A(n2955), .ZN(n3409) );
  AOI22_X1 U2606 ( .A1(datain[6]), .A2(n6009), .B1(n6571), .B2(
        \registers[22][6] ), .ZN(n2955) );
  INV_X1 U2607 ( .A(n2954), .ZN(n3410) );
  AOI22_X1 U2608 ( .A1(datain[7]), .A2(n6009), .B1(n6572), .B2(
        \registers[22][7] ), .ZN(n2954) );
  INV_X1 U2609 ( .A(n2953), .ZN(n3411) );
  AOI22_X1 U2610 ( .A1(datain[8]), .A2(n6009), .B1(n6572), .B2(
        \registers[22][8] ), .ZN(n2953) );
  INV_X1 U2611 ( .A(n2952), .ZN(n3412) );
  AOI22_X1 U2612 ( .A1(datain[9]), .A2(n6009), .B1(n6573), .B2(
        \registers[22][9] ), .ZN(n2952) );
  INV_X1 U2613 ( .A(n2951), .ZN(n3413) );
  AOI22_X1 U2614 ( .A1(datain[10]), .A2(n6009), .B1(n6573), .B2(
        \registers[22][10] ), .ZN(n2951) );
  INV_X1 U2615 ( .A(n2950), .ZN(n3414) );
  AOI22_X1 U2616 ( .A1(datain[11]), .A2(n6009), .B1(n6575), .B2(
        \registers[22][11] ), .ZN(n2950) );
  INV_X1 U2617 ( .A(n2949), .ZN(n3415) );
  AOI22_X1 U2618 ( .A1(datain[12]), .A2(n6010), .B1(n6569), .B2(
        \registers[22][12] ), .ZN(n2949) );
  INV_X1 U2619 ( .A(n2948), .ZN(n3416) );
  AOI22_X1 U2620 ( .A1(datain[13]), .A2(n6010), .B1(n6570), .B2(
        \registers[22][13] ), .ZN(n2948) );
  INV_X1 U2621 ( .A(n2947), .ZN(n3417) );
  AOI22_X1 U2622 ( .A1(datain[14]), .A2(n6010), .B1(n6571), .B2(
        \registers[22][14] ), .ZN(n2947) );
  INV_X1 U2623 ( .A(n2946), .ZN(n3418) );
  AOI22_X1 U2624 ( .A1(datain[15]), .A2(n6010), .B1(n6570), .B2(
        \registers[22][15] ), .ZN(n2946) );
  INV_X1 U2625 ( .A(n2945), .ZN(n3419) );
  AOI22_X1 U2626 ( .A1(datain[16]), .A2(n6010), .B1(n6572), .B2(
        \registers[22][16] ), .ZN(n2945) );
  INV_X1 U2627 ( .A(n2944), .ZN(n3420) );
  AOI22_X1 U2628 ( .A1(datain[17]), .A2(n6010), .B1(n6572), .B2(
        \registers[22][17] ), .ZN(n2944) );
  INV_X1 U2629 ( .A(n2943), .ZN(n3421) );
  AOI22_X1 U2630 ( .A1(datain[18]), .A2(n6010), .B1(n6573), .B2(
        \registers[22][18] ), .ZN(n2943) );
  INV_X1 U2631 ( .A(n2942), .ZN(n3422) );
  AOI22_X1 U2632 ( .A1(datain[19]), .A2(n6010), .B1(n6572), .B2(
        \registers[22][19] ), .ZN(n2942) );
  INV_X1 U2633 ( .A(n2941), .ZN(n3423) );
  AOI22_X1 U2634 ( .A1(datain[20]), .A2(n6010), .B1(n6574), .B2(
        \registers[22][20] ), .ZN(n2941) );
  INV_X1 U2635 ( .A(n2940), .ZN(n3424) );
  AOI22_X1 U2636 ( .A1(datain[21]), .A2(n6010), .B1(n6575), .B2(
        \registers[22][21] ), .ZN(n2940) );
  INV_X1 U2637 ( .A(n2939), .ZN(n3425) );
  AOI22_X1 U2638 ( .A1(datain[22]), .A2(n6010), .B1(n6574), .B2(
        \registers[22][22] ), .ZN(n2939) );
  INV_X1 U2639 ( .A(n2938), .ZN(n3426) );
  AOI22_X1 U2640 ( .A1(datain[23]), .A2(n6010), .B1(n6574), .B2(
        \registers[22][23] ), .ZN(n2938) );
  INV_X1 U2641 ( .A(n2937), .ZN(n3427) );
  AOI22_X1 U2642 ( .A1(datain[24]), .A2(n6011), .B1(n6575), .B2(
        \registers[22][24] ), .ZN(n2937) );
  INV_X1 U2643 ( .A(n2936), .ZN(n3428) );
  AOI22_X1 U2644 ( .A1(datain[25]), .A2(n6011), .B1(n6575), .B2(
        \registers[22][25] ), .ZN(n2936) );
  INV_X1 U2645 ( .A(n2935), .ZN(n3429) );
  AOI22_X1 U2646 ( .A1(datain[26]), .A2(n6011), .B1(n6569), .B2(
        \registers[22][26] ), .ZN(n2935) );
  INV_X1 U2647 ( .A(n2934), .ZN(n3430) );
  AOI22_X1 U2648 ( .A1(datain[27]), .A2(n6011), .B1(n6569), .B2(
        \registers[22][27] ), .ZN(n2934) );
  INV_X1 U2649 ( .A(n2933), .ZN(n3431) );
  AOI22_X1 U2650 ( .A1(datain[28]), .A2(n6011), .B1(n6569), .B2(
        \registers[22][28] ), .ZN(n2933) );
  INV_X1 U2651 ( .A(n2932), .ZN(n3432) );
  AOI22_X1 U2652 ( .A1(datain[29]), .A2(n6011), .B1(n6575), .B2(
        \registers[22][29] ), .ZN(n2932) );
  INV_X1 U2653 ( .A(n2931), .ZN(n3433) );
  AOI22_X1 U2654 ( .A1(datain[30]), .A2(n6011), .B1(n6570), .B2(
        \registers[22][30] ), .ZN(n2931) );
  INV_X1 U2655 ( .A(n2928), .ZN(n3434) );
  AOI22_X1 U2656 ( .A1(datain[31]), .A2(n6011), .B1(n6573), .B2(
        \registers[22][31] ), .ZN(n2928) );
  INV_X1 U2657 ( .A(n2927), .ZN(n3435) );
  AOI22_X1 U2658 ( .A1(datain[0]), .A2(n6012), .B1(n6578), .B2(
        \registers[21][0] ), .ZN(n2927) );
  INV_X1 U2659 ( .A(n2926), .ZN(n3436) );
  AOI22_X1 U2660 ( .A1(datain[1]), .A2(n6012), .B1(n6579), .B2(
        \registers[21][1] ), .ZN(n2926) );
  INV_X1 U2661 ( .A(n2925), .ZN(n3437) );
  AOI22_X1 U2662 ( .A1(datain[2]), .A2(n6012), .B1(n6580), .B2(
        \registers[21][2] ), .ZN(n2925) );
  INV_X1 U2663 ( .A(n2924), .ZN(n3438) );
  AOI22_X1 U2664 ( .A1(datain[3]), .A2(n6012), .B1(n6583), .B2(
        \registers[21][3] ), .ZN(n2924) );
  INV_X1 U2665 ( .A(n2923), .ZN(n3439) );
  AOI22_X1 U2666 ( .A1(datain[4]), .A2(n6012), .B1(n6579), .B2(
        \registers[21][4] ), .ZN(n2923) );
  INV_X1 U2667 ( .A(n2922), .ZN(n3440) );
  AOI22_X1 U2668 ( .A1(datain[5]), .A2(n6012), .B1(n6580), .B2(
        \registers[21][5] ), .ZN(n2922) );
  INV_X1 U2669 ( .A(n2921), .ZN(n3441) );
  AOI22_X1 U2670 ( .A1(datain[6]), .A2(n6012), .B1(n6580), .B2(
        \registers[21][6] ), .ZN(n2921) );
  INV_X1 U2671 ( .A(n2920), .ZN(n3442) );
  AOI22_X1 U2672 ( .A1(datain[7]), .A2(n6012), .B1(n6581), .B2(
        \registers[21][7] ), .ZN(n2920) );
  INV_X1 U2673 ( .A(n2919), .ZN(n3443) );
  AOI22_X1 U2674 ( .A1(datain[8]), .A2(n6012), .B1(n6581), .B2(
        \registers[21][8] ), .ZN(n2919) );
  INV_X1 U2675 ( .A(n2918), .ZN(n3444) );
  AOI22_X1 U2676 ( .A1(datain[9]), .A2(n6012), .B1(n6582), .B2(
        \registers[21][9] ), .ZN(n2918) );
  INV_X1 U2677 ( .A(n2917), .ZN(n3445) );
  AOI22_X1 U2678 ( .A1(datain[10]), .A2(n6012), .B1(n6582), .B2(
        \registers[21][10] ), .ZN(n2917) );
  INV_X1 U2679 ( .A(n2916), .ZN(n3446) );
  AOI22_X1 U2680 ( .A1(datain[11]), .A2(n6012), .B1(n6584), .B2(
        \registers[21][11] ), .ZN(n2916) );
  INV_X1 U2681 ( .A(n2915), .ZN(n3447) );
  AOI22_X1 U2682 ( .A1(datain[12]), .A2(n6013), .B1(n6578), .B2(
        \registers[21][12] ), .ZN(n2915) );
  INV_X1 U2683 ( .A(n2914), .ZN(n3448) );
  AOI22_X1 U2684 ( .A1(datain[13]), .A2(n6013), .B1(n6579), .B2(
        \registers[21][13] ), .ZN(n2914) );
  INV_X1 U2685 ( .A(n2913), .ZN(n3449) );
  AOI22_X1 U2686 ( .A1(datain[14]), .A2(n6013), .B1(n6580), .B2(
        \registers[21][14] ), .ZN(n2913) );
  INV_X1 U2687 ( .A(n2912), .ZN(n3450) );
  AOI22_X1 U2688 ( .A1(datain[15]), .A2(n6013), .B1(n6579), .B2(
        \registers[21][15] ), .ZN(n2912) );
  INV_X1 U2689 ( .A(n2911), .ZN(n3451) );
  AOI22_X1 U2690 ( .A1(datain[16]), .A2(n6013), .B1(n6581), .B2(
        \registers[21][16] ), .ZN(n2911) );
  INV_X1 U2691 ( .A(n2910), .ZN(n3452) );
  AOI22_X1 U2692 ( .A1(datain[17]), .A2(n6013), .B1(n6581), .B2(
        \registers[21][17] ), .ZN(n2910) );
  INV_X1 U2693 ( .A(n2909), .ZN(n3453) );
  AOI22_X1 U2694 ( .A1(datain[18]), .A2(n6013), .B1(n6582), .B2(
        \registers[21][18] ), .ZN(n2909) );
  INV_X1 U2695 ( .A(n2908), .ZN(n3454) );
  AOI22_X1 U2696 ( .A1(datain[19]), .A2(n6013), .B1(n6581), .B2(
        \registers[21][19] ), .ZN(n2908) );
  INV_X1 U2697 ( .A(n2907), .ZN(n3455) );
  AOI22_X1 U2698 ( .A1(datain[20]), .A2(n6013), .B1(n6583), .B2(
        \registers[21][20] ), .ZN(n2907) );
  INV_X1 U2699 ( .A(n2906), .ZN(n3456) );
  AOI22_X1 U2700 ( .A1(datain[21]), .A2(n6013), .B1(n6584), .B2(
        \registers[21][21] ), .ZN(n2906) );
  INV_X1 U2701 ( .A(n2905), .ZN(n3457) );
  AOI22_X1 U2702 ( .A1(datain[22]), .A2(n6013), .B1(n6583), .B2(
        \registers[21][22] ), .ZN(n2905) );
  INV_X1 U2703 ( .A(n2904), .ZN(n3458) );
  AOI22_X1 U2704 ( .A1(datain[23]), .A2(n6013), .B1(n6583), .B2(
        \registers[21][23] ), .ZN(n2904) );
  INV_X1 U2705 ( .A(n2903), .ZN(n3459) );
  AOI22_X1 U2706 ( .A1(datain[24]), .A2(n6014), .B1(n6584), .B2(
        \registers[21][24] ), .ZN(n2903) );
  INV_X1 U2707 ( .A(n2902), .ZN(n3460) );
  AOI22_X1 U2708 ( .A1(datain[25]), .A2(n6014), .B1(n6584), .B2(
        \registers[21][25] ), .ZN(n2902) );
  INV_X1 U2709 ( .A(n2901), .ZN(n3461) );
  AOI22_X1 U2710 ( .A1(datain[26]), .A2(n6014), .B1(n6578), .B2(
        \registers[21][26] ), .ZN(n2901) );
  INV_X1 U2711 ( .A(n2900), .ZN(n3462) );
  AOI22_X1 U2712 ( .A1(datain[27]), .A2(n6014), .B1(n6578), .B2(
        \registers[21][27] ), .ZN(n2900) );
  INV_X1 U2713 ( .A(n2899), .ZN(n3463) );
  AOI22_X1 U2714 ( .A1(datain[28]), .A2(n6014), .B1(n6578), .B2(
        \registers[21][28] ), .ZN(n2899) );
  INV_X1 U2715 ( .A(n2898), .ZN(n3464) );
  AOI22_X1 U2716 ( .A1(datain[29]), .A2(n6014), .B1(n6584), .B2(
        \registers[21][29] ), .ZN(n2898) );
  INV_X1 U2717 ( .A(n2897), .ZN(n3465) );
  AOI22_X1 U2718 ( .A1(datain[30]), .A2(n6014), .B1(n6579), .B2(
        \registers[21][30] ), .ZN(n2897) );
  INV_X1 U2719 ( .A(n2894), .ZN(n3466) );
  AOI22_X1 U2720 ( .A1(datain[31]), .A2(n6014), .B1(n6582), .B2(
        \registers[21][31] ), .ZN(n2894) );
  INV_X1 U2721 ( .A(n2892), .ZN(n3467) );
  AOI22_X1 U2722 ( .A1(datain[0]), .A2(n6015), .B1(n6587), .B2(
        \registers[20][0] ), .ZN(n2892) );
  INV_X1 U2723 ( .A(n2891), .ZN(n3468) );
  AOI22_X1 U2724 ( .A1(datain[1]), .A2(n6015), .B1(n6588), .B2(
        \registers[20][1] ), .ZN(n2891) );
  INV_X1 U2725 ( .A(n2890), .ZN(n3469) );
  AOI22_X1 U2726 ( .A1(datain[2]), .A2(n6015), .B1(n6589), .B2(
        \registers[20][2] ), .ZN(n2890) );
  INV_X1 U2727 ( .A(n2889), .ZN(n3470) );
  AOI22_X1 U2728 ( .A1(datain[3]), .A2(n6015), .B1(n6592), .B2(
        \registers[20][3] ), .ZN(n2889) );
  INV_X1 U2729 ( .A(n2888), .ZN(n3471) );
  AOI22_X1 U2730 ( .A1(datain[4]), .A2(n6015), .B1(n6588), .B2(
        \registers[20][4] ), .ZN(n2888) );
  INV_X1 U2731 ( .A(n2887), .ZN(n3472) );
  AOI22_X1 U2732 ( .A1(datain[5]), .A2(n6015), .B1(n6589), .B2(
        \registers[20][5] ), .ZN(n2887) );
  INV_X1 U2733 ( .A(n2886), .ZN(n3473) );
  AOI22_X1 U2734 ( .A1(datain[6]), .A2(n6015), .B1(n6589), .B2(
        \registers[20][6] ), .ZN(n2886) );
  INV_X1 U2735 ( .A(n2885), .ZN(n3474) );
  AOI22_X1 U2736 ( .A1(datain[7]), .A2(n6015), .B1(n6590), .B2(
        \registers[20][7] ), .ZN(n2885) );
  INV_X1 U2737 ( .A(n2884), .ZN(n3475) );
  AOI22_X1 U2738 ( .A1(datain[8]), .A2(n6015), .B1(n6590), .B2(
        \registers[20][8] ), .ZN(n2884) );
  INV_X1 U2739 ( .A(n2883), .ZN(n3476) );
  AOI22_X1 U2740 ( .A1(datain[9]), .A2(n6015), .B1(n6591), .B2(
        \registers[20][9] ), .ZN(n2883) );
  INV_X1 U2741 ( .A(n2882), .ZN(n3477) );
  AOI22_X1 U2742 ( .A1(datain[10]), .A2(n6015), .B1(n6591), .B2(
        \registers[20][10] ), .ZN(n2882) );
  INV_X1 U2743 ( .A(n2881), .ZN(n3478) );
  AOI22_X1 U2744 ( .A1(datain[11]), .A2(n6015), .B1(n6593), .B2(
        \registers[20][11] ), .ZN(n2881) );
  INV_X1 U2745 ( .A(n2880), .ZN(n3479) );
  AOI22_X1 U2746 ( .A1(datain[12]), .A2(n6016), .B1(n6587), .B2(
        \registers[20][12] ), .ZN(n2880) );
  INV_X1 U2747 ( .A(n2879), .ZN(n3480) );
  AOI22_X1 U2748 ( .A1(datain[13]), .A2(n6016), .B1(n6588), .B2(
        \registers[20][13] ), .ZN(n2879) );
  INV_X1 U2749 ( .A(n2878), .ZN(n3481) );
  AOI22_X1 U2750 ( .A1(datain[14]), .A2(n6016), .B1(n6589), .B2(
        \registers[20][14] ), .ZN(n2878) );
  INV_X1 U2751 ( .A(n2877), .ZN(n3482) );
  AOI22_X1 U2752 ( .A1(datain[15]), .A2(n6016), .B1(n6588), .B2(
        \registers[20][15] ), .ZN(n2877) );
  INV_X1 U2753 ( .A(n2876), .ZN(n3483) );
  AOI22_X1 U2754 ( .A1(datain[16]), .A2(n6016), .B1(n6590), .B2(
        \registers[20][16] ), .ZN(n2876) );
  INV_X1 U2755 ( .A(n2875), .ZN(n3484) );
  AOI22_X1 U2756 ( .A1(datain[17]), .A2(n6016), .B1(n6590), .B2(
        \registers[20][17] ), .ZN(n2875) );
  INV_X1 U2757 ( .A(n2874), .ZN(n3485) );
  AOI22_X1 U2758 ( .A1(datain[18]), .A2(n6016), .B1(n6591), .B2(
        \registers[20][18] ), .ZN(n2874) );
  INV_X1 U2759 ( .A(n2873), .ZN(n3486) );
  AOI22_X1 U2760 ( .A1(datain[19]), .A2(n6016), .B1(n6590), .B2(
        \registers[20][19] ), .ZN(n2873) );
  INV_X1 U2761 ( .A(n2872), .ZN(n3487) );
  AOI22_X1 U2762 ( .A1(datain[20]), .A2(n6016), .B1(n6592), .B2(
        \registers[20][20] ), .ZN(n2872) );
  INV_X1 U2763 ( .A(n2871), .ZN(n3488) );
  AOI22_X1 U2764 ( .A1(datain[21]), .A2(n6016), .B1(n6593), .B2(
        \registers[20][21] ), .ZN(n2871) );
  INV_X1 U2765 ( .A(n2870), .ZN(n3489) );
  AOI22_X1 U2766 ( .A1(datain[22]), .A2(n6016), .B1(n6592), .B2(
        \registers[20][22] ), .ZN(n2870) );
  INV_X1 U2767 ( .A(n2869), .ZN(n3490) );
  AOI22_X1 U2768 ( .A1(datain[23]), .A2(n6016), .B1(n6592), .B2(
        \registers[20][23] ), .ZN(n2869) );
  INV_X1 U2769 ( .A(n2868), .ZN(n3491) );
  AOI22_X1 U2770 ( .A1(datain[24]), .A2(n6017), .B1(n6593), .B2(
        \registers[20][24] ), .ZN(n2868) );
  INV_X1 U2771 ( .A(n2867), .ZN(n3492) );
  AOI22_X1 U2772 ( .A1(datain[25]), .A2(n6017), .B1(n6593), .B2(
        \registers[20][25] ), .ZN(n2867) );
  INV_X1 U2773 ( .A(n2866), .ZN(n3493) );
  AOI22_X1 U2774 ( .A1(datain[26]), .A2(n6017), .B1(n6587), .B2(
        \registers[20][26] ), .ZN(n2866) );
  INV_X1 U2775 ( .A(n2865), .ZN(n3494) );
  AOI22_X1 U2776 ( .A1(datain[27]), .A2(n6017), .B1(n6587), .B2(
        \registers[20][27] ), .ZN(n2865) );
  INV_X1 U2777 ( .A(n2864), .ZN(n3495) );
  AOI22_X1 U2778 ( .A1(datain[28]), .A2(n6017), .B1(n6587), .B2(
        \registers[20][28] ), .ZN(n2864) );
  INV_X1 U2779 ( .A(n2863), .ZN(n3496) );
  AOI22_X1 U2780 ( .A1(datain[29]), .A2(n6017), .B1(n6593), .B2(
        \registers[20][29] ), .ZN(n2863) );
  INV_X1 U2781 ( .A(n2862), .ZN(n3497) );
  AOI22_X1 U2782 ( .A1(datain[30]), .A2(n6017), .B1(n6588), .B2(
        \registers[20][30] ), .ZN(n2862) );
  INV_X1 U2783 ( .A(n2859), .ZN(n3498) );
  AOI22_X1 U2784 ( .A1(datain[31]), .A2(n6017), .B1(n6591), .B2(
        \registers[20][31] ), .ZN(n2859) );
  INV_X1 U2785 ( .A(n2718), .ZN(n3627) );
  AOI22_X1 U2786 ( .A1(datain[0]), .A2(n6030), .B1(n6629), .B2(
        \registers[15][0] ), .ZN(n2718) );
  INV_X1 U2787 ( .A(n2717), .ZN(n3628) );
  AOI22_X1 U2788 ( .A1(datain[1]), .A2(n6030), .B1(n6630), .B2(
        \registers[15][1] ), .ZN(n2717) );
  INV_X1 U2789 ( .A(n2716), .ZN(n3629) );
  AOI22_X1 U2790 ( .A1(datain[2]), .A2(n6030), .B1(n6631), .B2(
        \registers[15][2] ), .ZN(n2716) );
  INV_X1 U2791 ( .A(n2715), .ZN(n3630) );
  AOI22_X1 U2792 ( .A1(datain[3]), .A2(n6030), .B1(n6634), .B2(
        \registers[15][3] ), .ZN(n2715) );
  INV_X1 U2793 ( .A(n2714), .ZN(n3631) );
  AOI22_X1 U2794 ( .A1(datain[4]), .A2(n6030), .B1(n6630), .B2(
        \registers[15][4] ), .ZN(n2714) );
  INV_X1 U2795 ( .A(n2713), .ZN(n3632) );
  AOI22_X1 U2796 ( .A1(datain[5]), .A2(n6030), .B1(n6631), .B2(
        \registers[15][5] ), .ZN(n2713) );
  INV_X1 U2797 ( .A(n2712), .ZN(n3633) );
  AOI22_X1 U2798 ( .A1(datain[6]), .A2(n6030), .B1(n6631), .B2(
        \registers[15][6] ), .ZN(n2712) );
  INV_X1 U2799 ( .A(n2711), .ZN(n3634) );
  AOI22_X1 U2800 ( .A1(datain[7]), .A2(n6030), .B1(n6632), .B2(
        \registers[15][7] ), .ZN(n2711) );
  INV_X1 U2801 ( .A(n2710), .ZN(n3635) );
  AOI22_X1 U2802 ( .A1(datain[8]), .A2(n6030), .B1(n6632), .B2(
        \registers[15][8] ), .ZN(n2710) );
  INV_X1 U2803 ( .A(n2709), .ZN(n3636) );
  AOI22_X1 U2804 ( .A1(datain[9]), .A2(n6030), .B1(n6633), .B2(
        \registers[15][9] ), .ZN(n2709) );
  INV_X1 U2805 ( .A(n2708), .ZN(n3637) );
  AOI22_X1 U2806 ( .A1(datain[10]), .A2(n6030), .B1(n6633), .B2(
        \registers[15][10] ), .ZN(n2708) );
  INV_X1 U2807 ( .A(n2707), .ZN(n3638) );
  AOI22_X1 U2808 ( .A1(datain[11]), .A2(n6030), .B1(n6635), .B2(
        \registers[15][11] ), .ZN(n2707) );
  INV_X1 U2809 ( .A(n2706), .ZN(n3639) );
  AOI22_X1 U2810 ( .A1(datain[12]), .A2(n6031), .B1(n6629), .B2(
        \registers[15][12] ), .ZN(n2706) );
  INV_X1 U2811 ( .A(n2705), .ZN(n3640) );
  AOI22_X1 U2812 ( .A1(datain[13]), .A2(n6031), .B1(n6630), .B2(
        \registers[15][13] ), .ZN(n2705) );
  INV_X1 U2813 ( .A(n2704), .ZN(n3641) );
  AOI22_X1 U2814 ( .A1(datain[14]), .A2(n6031), .B1(n6631), .B2(
        \registers[15][14] ), .ZN(n2704) );
  INV_X1 U2815 ( .A(n2703), .ZN(n3642) );
  AOI22_X1 U2816 ( .A1(datain[15]), .A2(n6031), .B1(n6630), .B2(
        \registers[15][15] ), .ZN(n2703) );
  INV_X1 U2817 ( .A(n2702), .ZN(n3643) );
  AOI22_X1 U2818 ( .A1(datain[16]), .A2(n6031), .B1(n6632), .B2(
        \registers[15][16] ), .ZN(n2702) );
  INV_X1 U2819 ( .A(n2701), .ZN(n3644) );
  AOI22_X1 U2820 ( .A1(datain[17]), .A2(n6031), .B1(n6632), .B2(
        \registers[15][17] ), .ZN(n2701) );
  INV_X1 U2821 ( .A(n2700), .ZN(n3645) );
  AOI22_X1 U2822 ( .A1(datain[18]), .A2(n6031), .B1(n6633), .B2(
        \registers[15][18] ), .ZN(n2700) );
  INV_X1 U2823 ( .A(n2699), .ZN(n3646) );
  AOI22_X1 U2824 ( .A1(datain[19]), .A2(n6031), .B1(n6632), .B2(
        \registers[15][19] ), .ZN(n2699) );
  INV_X1 U2825 ( .A(n2698), .ZN(n3647) );
  AOI22_X1 U2826 ( .A1(datain[20]), .A2(n6031), .B1(n6634), .B2(
        \registers[15][20] ), .ZN(n2698) );
  INV_X1 U2827 ( .A(n2697), .ZN(n3648) );
  AOI22_X1 U2828 ( .A1(datain[21]), .A2(n6031), .B1(n6635), .B2(
        \registers[15][21] ), .ZN(n2697) );
  INV_X1 U2829 ( .A(n2696), .ZN(n3649) );
  AOI22_X1 U2830 ( .A1(datain[22]), .A2(n6031), .B1(n6634), .B2(
        \registers[15][22] ), .ZN(n2696) );
  INV_X1 U2831 ( .A(n2695), .ZN(n3650) );
  AOI22_X1 U2832 ( .A1(datain[23]), .A2(n6031), .B1(n6634), .B2(
        \registers[15][23] ), .ZN(n2695) );
  INV_X1 U2833 ( .A(n2694), .ZN(n3651) );
  AOI22_X1 U2834 ( .A1(datain[24]), .A2(n6032), .B1(n6635), .B2(
        \registers[15][24] ), .ZN(n2694) );
  INV_X1 U2835 ( .A(n2693), .ZN(n3652) );
  AOI22_X1 U2836 ( .A1(datain[25]), .A2(n6032), .B1(n6635), .B2(
        \registers[15][25] ), .ZN(n2693) );
  INV_X1 U2837 ( .A(n2692), .ZN(n3653) );
  AOI22_X1 U2838 ( .A1(datain[26]), .A2(n6032), .B1(n6629), .B2(
        \registers[15][26] ), .ZN(n2692) );
  INV_X1 U2839 ( .A(n2691), .ZN(n3654) );
  AOI22_X1 U2840 ( .A1(datain[27]), .A2(n6032), .B1(n6629), .B2(
        \registers[15][27] ), .ZN(n2691) );
  INV_X1 U2841 ( .A(n2690), .ZN(n3655) );
  AOI22_X1 U2842 ( .A1(datain[28]), .A2(n6032), .B1(n6629), .B2(
        \registers[15][28] ), .ZN(n2690) );
  INV_X1 U2843 ( .A(n2689), .ZN(n3656) );
  AOI22_X1 U2844 ( .A1(datain[29]), .A2(n6032), .B1(n6635), .B2(
        \registers[15][29] ), .ZN(n2689) );
  INV_X1 U2845 ( .A(n2688), .ZN(n3657) );
  AOI22_X1 U2846 ( .A1(datain[30]), .A2(n6032), .B1(n6630), .B2(
        \registers[15][30] ), .ZN(n2688) );
  INV_X1 U2847 ( .A(n2685), .ZN(n3658) );
  AOI22_X1 U2848 ( .A1(datain[31]), .A2(n6032), .B1(n6633), .B2(
        \registers[15][31] ), .ZN(n2685) );
  INV_X1 U2849 ( .A(n2684), .ZN(n3659) );
  AOI22_X1 U2850 ( .A1(datain[0]), .A2(n6033), .B1(n6638), .B2(
        \registers[14][0] ), .ZN(n2684) );
  INV_X1 U2851 ( .A(n2683), .ZN(n3660) );
  AOI22_X1 U2852 ( .A1(datain[1]), .A2(n6033), .B1(n6639), .B2(
        \registers[14][1] ), .ZN(n2683) );
  INV_X1 U2853 ( .A(n2682), .ZN(n3661) );
  AOI22_X1 U2854 ( .A1(datain[2]), .A2(n6033), .B1(n6640), .B2(
        \registers[14][2] ), .ZN(n2682) );
  INV_X1 U2855 ( .A(n2681), .ZN(n3662) );
  AOI22_X1 U2856 ( .A1(datain[3]), .A2(n6033), .B1(n6643), .B2(
        \registers[14][3] ), .ZN(n2681) );
  INV_X1 U2857 ( .A(n2680), .ZN(n3663) );
  AOI22_X1 U2858 ( .A1(datain[4]), .A2(n6033), .B1(n6639), .B2(
        \registers[14][4] ), .ZN(n2680) );
  INV_X1 U2859 ( .A(n2679), .ZN(n3664) );
  AOI22_X1 U2860 ( .A1(datain[5]), .A2(n6033), .B1(n6640), .B2(
        \registers[14][5] ), .ZN(n2679) );
  INV_X1 U2861 ( .A(n2678), .ZN(n3665) );
  AOI22_X1 U2862 ( .A1(datain[6]), .A2(n6033), .B1(n6640), .B2(
        \registers[14][6] ), .ZN(n2678) );
  INV_X1 U2863 ( .A(n2677), .ZN(n3666) );
  AOI22_X1 U2864 ( .A1(datain[7]), .A2(n6033), .B1(n6641), .B2(
        \registers[14][7] ), .ZN(n2677) );
  INV_X1 U2865 ( .A(n2676), .ZN(n3667) );
  AOI22_X1 U2866 ( .A1(datain[8]), .A2(n6033), .B1(n6641), .B2(
        \registers[14][8] ), .ZN(n2676) );
  INV_X1 U2867 ( .A(n2675), .ZN(n3668) );
  AOI22_X1 U2868 ( .A1(datain[9]), .A2(n6033), .B1(n6642), .B2(
        \registers[14][9] ), .ZN(n2675) );
  INV_X1 U2869 ( .A(n2674), .ZN(n3669) );
  AOI22_X1 U2870 ( .A1(datain[10]), .A2(n6033), .B1(n6642), .B2(
        \registers[14][10] ), .ZN(n2674) );
  INV_X1 U2871 ( .A(n2673), .ZN(n3670) );
  AOI22_X1 U2872 ( .A1(datain[11]), .A2(n6033), .B1(n6644), .B2(
        \registers[14][11] ), .ZN(n2673) );
  INV_X1 U2873 ( .A(n2672), .ZN(n3671) );
  AOI22_X1 U2874 ( .A1(datain[12]), .A2(n6034), .B1(n6638), .B2(
        \registers[14][12] ), .ZN(n2672) );
  INV_X1 U2875 ( .A(n2671), .ZN(n3672) );
  AOI22_X1 U2876 ( .A1(datain[13]), .A2(n6034), .B1(n6639), .B2(
        \registers[14][13] ), .ZN(n2671) );
  INV_X1 U2877 ( .A(n2670), .ZN(n3673) );
  AOI22_X1 U2878 ( .A1(datain[14]), .A2(n6034), .B1(n6640), .B2(
        \registers[14][14] ), .ZN(n2670) );
  INV_X1 U2879 ( .A(n2669), .ZN(n3674) );
  AOI22_X1 U2880 ( .A1(datain[15]), .A2(n6034), .B1(n6639), .B2(
        \registers[14][15] ), .ZN(n2669) );
  INV_X1 U2881 ( .A(n2668), .ZN(n3675) );
  AOI22_X1 U2882 ( .A1(datain[16]), .A2(n6034), .B1(n6641), .B2(
        \registers[14][16] ), .ZN(n2668) );
  INV_X1 U2883 ( .A(n2667), .ZN(n3676) );
  AOI22_X1 U2884 ( .A1(datain[17]), .A2(n6034), .B1(n6641), .B2(
        \registers[14][17] ), .ZN(n2667) );
  INV_X1 U2885 ( .A(n2666), .ZN(n3677) );
  AOI22_X1 U2886 ( .A1(datain[18]), .A2(n6034), .B1(n6642), .B2(
        \registers[14][18] ), .ZN(n2666) );
  INV_X1 U2887 ( .A(n2665), .ZN(n3678) );
  AOI22_X1 U2888 ( .A1(datain[19]), .A2(n6034), .B1(n6641), .B2(
        \registers[14][19] ), .ZN(n2665) );
  INV_X1 U2889 ( .A(n2664), .ZN(n3679) );
  AOI22_X1 U2890 ( .A1(datain[20]), .A2(n6034), .B1(n6643), .B2(
        \registers[14][20] ), .ZN(n2664) );
  INV_X1 U2891 ( .A(n2663), .ZN(n3680) );
  AOI22_X1 U2892 ( .A1(datain[21]), .A2(n6034), .B1(n6644), .B2(
        \registers[14][21] ), .ZN(n2663) );
  INV_X1 U2893 ( .A(n2662), .ZN(n3681) );
  AOI22_X1 U2894 ( .A1(datain[22]), .A2(n6034), .B1(n6643), .B2(
        \registers[14][22] ), .ZN(n2662) );
  INV_X1 U2895 ( .A(n2661), .ZN(n3682) );
  AOI22_X1 U2896 ( .A1(datain[23]), .A2(n6034), .B1(n6643), .B2(
        \registers[14][23] ), .ZN(n2661) );
  INV_X1 U2897 ( .A(n2660), .ZN(n3683) );
  AOI22_X1 U2898 ( .A1(datain[24]), .A2(n6035), .B1(n6644), .B2(
        \registers[14][24] ), .ZN(n2660) );
  INV_X1 U2899 ( .A(n2659), .ZN(n3684) );
  AOI22_X1 U2900 ( .A1(datain[25]), .A2(n6035), .B1(n6644), .B2(
        \registers[14][25] ), .ZN(n2659) );
  INV_X1 U2901 ( .A(n2658), .ZN(n3685) );
  AOI22_X1 U2902 ( .A1(datain[26]), .A2(n6035), .B1(n6638), .B2(
        \registers[14][26] ), .ZN(n2658) );
  INV_X1 U2903 ( .A(n2657), .ZN(n3686) );
  AOI22_X1 U2904 ( .A1(datain[27]), .A2(n6035), .B1(n6638), .B2(
        \registers[14][27] ), .ZN(n2657) );
  INV_X1 U2905 ( .A(n2656), .ZN(n3687) );
  AOI22_X1 U2906 ( .A1(datain[28]), .A2(n6035), .B1(n6638), .B2(
        \registers[14][28] ), .ZN(n2656) );
  INV_X1 U2907 ( .A(n2655), .ZN(n3688) );
  AOI22_X1 U2908 ( .A1(datain[29]), .A2(n6035), .B1(n6644), .B2(
        \registers[14][29] ), .ZN(n2655) );
  INV_X1 U2909 ( .A(n2654), .ZN(n3689) );
  AOI22_X1 U2910 ( .A1(datain[30]), .A2(n6035), .B1(n6639), .B2(
        \registers[14][30] ), .ZN(n2654) );
  INV_X1 U2911 ( .A(n2651), .ZN(n3690) );
  AOI22_X1 U2912 ( .A1(datain[31]), .A2(n6035), .B1(n6642), .B2(
        \registers[14][31] ), .ZN(n2651) );
  INV_X1 U2913 ( .A(n2650), .ZN(n3691) );
  AOI22_X1 U2914 ( .A1(datain[0]), .A2(n6036), .B1(n6647), .B2(
        \registers[13][0] ), .ZN(n2650) );
  INV_X1 U2915 ( .A(n2649), .ZN(n3692) );
  AOI22_X1 U2916 ( .A1(datain[1]), .A2(n6036), .B1(n6648), .B2(
        \registers[13][1] ), .ZN(n2649) );
  INV_X1 U2917 ( .A(n2648), .ZN(n3693) );
  AOI22_X1 U2918 ( .A1(datain[2]), .A2(n6036), .B1(n6649), .B2(
        \registers[13][2] ), .ZN(n2648) );
  INV_X1 U2919 ( .A(n2647), .ZN(n3694) );
  AOI22_X1 U2920 ( .A1(datain[3]), .A2(n6036), .B1(n6652), .B2(
        \registers[13][3] ), .ZN(n2647) );
  INV_X1 U2921 ( .A(n2646), .ZN(n3695) );
  AOI22_X1 U2922 ( .A1(datain[4]), .A2(n6036), .B1(n6648), .B2(
        \registers[13][4] ), .ZN(n2646) );
  INV_X1 U2923 ( .A(n2645), .ZN(n3696) );
  AOI22_X1 U2924 ( .A1(datain[5]), .A2(n6036), .B1(n6649), .B2(
        \registers[13][5] ), .ZN(n2645) );
  INV_X1 U2925 ( .A(n2644), .ZN(n3697) );
  AOI22_X1 U2926 ( .A1(datain[6]), .A2(n6036), .B1(n6649), .B2(
        \registers[13][6] ), .ZN(n2644) );
  INV_X1 U2927 ( .A(n2643), .ZN(n3698) );
  AOI22_X1 U2928 ( .A1(datain[7]), .A2(n6036), .B1(n6650), .B2(
        \registers[13][7] ), .ZN(n2643) );
  INV_X1 U2929 ( .A(n2642), .ZN(n3699) );
  AOI22_X1 U2930 ( .A1(datain[8]), .A2(n6036), .B1(n6650), .B2(
        \registers[13][8] ), .ZN(n2642) );
  INV_X1 U2931 ( .A(n2641), .ZN(n3700) );
  AOI22_X1 U2932 ( .A1(datain[9]), .A2(n6036), .B1(n6651), .B2(
        \registers[13][9] ), .ZN(n2641) );
  INV_X1 U2933 ( .A(n2640), .ZN(n3701) );
  AOI22_X1 U2934 ( .A1(datain[10]), .A2(n6036), .B1(n6651), .B2(
        \registers[13][10] ), .ZN(n2640) );
  INV_X1 U2935 ( .A(n2639), .ZN(n3702) );
  AOI22_X1 U2936 ( .A1(datain[11]), .A2(n6036), .B1(n6653), .B2(
        \registers[13][11] ), .ZN(n2639) );
  INV_X1 U2937 ( .A(n2638), .ZN(n3703) );
  AOI22_X1 U2938 ( .A1(datain[12]), .A2(n6037), .B1(n6647), .B2(
        \registers[13][12] ), .ZN(n2638) );
  INV_X1 U2939 ( .A(n2637), .ZN(n3704) );
  AOI22_X1 U2940 ( .A1(datain[13]), .A2(n6037), .B1(n6648), .B2(
        \registers[13][13] ), .ZN(n2637) );
  INV_X1 U2941 ( .A(n2636), .ZN(n3705) );
  AOI22_X1 U2942 ( .A1(datain[14]), .A2(n6037), .B1(n6649), .B2(
        \registers[13][14] ), .ZN(n2636) );
  INV_X1 U2943 ( .A(n2635), .ZN(n3706) );
  AOI22_X1 U2944 ( .A1(datain[15]), .A2(n6037), .B1(n6648), .B2(
        \registers[13][15] ), .ZN(n2635) );
  INV_X1 U2945 ( .A(n2634), .ZN(n3707) );
  AOI22_X1 U2946 ( .A1(datain[16]), .A2(n6037), .B1(n6650), .B2(
        \registers[13][16] ), .ZN(n2634) );
  INV_X1 U2947 ( .A(n2633), .ZN(n3708) );
  AOI22_X1 U2948 ( .A1(datain[17]), .A2(n6037), .B1(n6650), .B2(
        \registers[13][17] ), .ZN(n2633) );
  INV_X1 U2949 ( .A(n2632), .ZN(n3709) );
  AOI22_X1 U2950 ( .A1(datain[18]), .A2(n6037), .B1(n6651), .B2(
        \registers[13][18] ), .ZN(n2632) );
  INV_X1 U2951 ( .A(n2631), .ZN(n3710) );
  AOI22_X1 U2952 ( .A1(datain[19]), .A2(n6037), .B1(n6650), .B2(
        \registers[13][19] ), .ZN(n2631) );
  INV_X1 U2953 ( .A(n2630), .ZN(n3711) );
  AOI22_X1 U2954 ( .A1(datain[20]), .A2(n6037), .B1(n6652), .B2(
        \registers[13][20] ), .ZN(n2630) );
  INV_X1 U2955 ( .A(n2629), .ZN(n3712) );
  AOI22_X1 U2956 ( .A1(datain[21]), .A2(n6037), .B1(n6653), .B2(
        \registers[13][21] ), .ZN(n2629) );
  INV_X1 U2957 ( .A(n2628), .ZN(n3713) );
  AOI22_X1 U2958 ( .A1(datain[22]), .A2(n6037), .B1(n6652), .B2(
        \registers[13][22] ), .ZN(n2628) );
  INV_X1 U2959 ( .A(n2627), .ZN(n3714) );
  AOI22_X1 U2960 ( .A1(datain[23]), .A2(n6037), .B1(n6652), .B2(
        \registers[13][23] ), .ZN(n2627) );
  INV_X1 U2961 ( .A(n2626), .ZN(n3715) );
  AOI22_X1 U2962 ( .A1(datain[24]), .A2(n6038), .B1(n6653), .B2(
        \registers[13][24] ), .ZN(n2626) );
  INV_X1 U2963 ( .A(n2625), .ZN(n3716) );
  AOI22_X1 U2964 ( .A1(datain[25]), .A2(n6038), .B1(n6653), .B2(
        \registers[13][25] ), .ZN(n2625) );
  INV_X1 U2965 ( .A(n2624), .ZN(n3717) );
  AOI22_X1 U2966 ( .A1(datain[26]), .A2(n6038), .B1(n6647), .B2(
        \registers[13][26] ), .ZN(n2624) );
  INV_X1 U2967 ( .A(n2623), .ZN(n3718) );
  AOI22_X1 U2968 ( .A1(datain[27]), .A2(n6038), .B1(n6647), .B2(
        \registers[13][27] ), .ZN(n2623) );
  INV_X1 U2969 ( .A(n2622), .ZN(n3719) );
  AOI22_X1 U2970 ( .A1(datain[28]), .A2(n6038), .B1(n6647), .B2(
        \registers[13][28] ), .ZN(n2622) );
  INV_X1 U2971 ( .A(n2621), .ZN(n3720) );
  AOI22_X1 U2972 ( .A1(datain[29]), .A2(n6038), .B1(n6653), .B2(
        \registers[13][29] ), .ZN(n2621) );
  INV_X1 U2973 ( .A(n2620), .ZN(n3721) );
  AOI22_X1 U2974 ( .A1(datain[30]), .A2(n6038), .B1(n6648), .B2(
        \registers[13][30] ), .ZN(n2620) );
  INV_X1 U2975 ( .A(n2617), .ZN(n3722) );
  AOI22_X1 U2976 ( .A1(datain[31]), .A2(n6038), .B1(n6651), .B2(
        \registers[13][31] ), .ZN(n2617) );
  INV_X1 U2977 ( .A(n2615), .ZN(n3723) );
  AOI22_X1 U2978 ( .A1(datain[0]), .A2(n6039), .B1(n6656), .B2(
        \registers[12][0] ), .ZN(n2615) );
  INV_X1 U2979 ( .A(n2614), .ZN(n3724) );
  AOI22_X1 U2980 ( .A1(datain[1]), .A2(n6039), .B1(n6657), .B2(
        \registers[12][1] ), .ZN(n2614) );
  INV_X1 U2981 ( .A(n2613), .ZN(n3725) );
  AOI22_X1 U2982 ( .A1(datain[2]), .A2(n6039), .B1(n6658), .B2(
        \registers[12][2] ), .ZN(n2613) );
  INV_X1 U2983 ( .A(n2612), .ZN(n3726) );
  AOI22_X1 U2984 ( .A1(datain[3]), .A2(n6039), .B1(n6661), .B2(
        \registers[12][3] ), .ZN(n2612) );
  INV_X1 U2985 ( .A(n2611), .ZN(n3727) );
  AOI22_X1 U2986 ( .A1(datain[4]), .A2(n6039), .B1(n6657), .B2(
        \registers[12][4] ), .ZN(n2611) );
  INV_X1 U2987 ( .A(n2610), .ZN(n3728) );
  AOI22_X1 U2988 ( .A1(datain[5]), .A2(n6039), .B1(n6658), .B2(
        \registers[12][5] ), .ZN(n2610) );
  INV_X1 U2989 ( .A(n2609), .ZN(n3729) );
  AOI22_X1 U2990 ( .A1(datain[6]), .A2(n6039), .B1(n6658), .B2(
        \registers[12][6] ), .ZN(n2609) );
  INV_X1 U2991 ( .A(n2608), .ZN(n3730) );
  AOI22_X1 U2992 ( .A1(datain[7]), .A2(n6039), .B1(n6659), .B2(
        \registers[12][7] ), .ZN(n2608) );
  INV_X1 U2993 ( .A(n2607), .ZN(n3731) );
  AOI22_X1 U2994 ( .A1(datain[8]), .A2(n6039), .B1(n6659), .B2(
        \registers[12][8] ), .ZN(n2607) );
  INV_X1 U2995 ( .A(n2606), .ZN(n3732) );
  AOI22_X1 U2996 ( .A1(datain[9]), .A2(n6039), .B1(n6660), .B2(
        \registers[12][9] ), .ZN(n2606) );
  INV_X1 U2997 ( .A(n2605), .ZN(n3733) );
  AOI22_X1 U2998 ( .A1(datain[10]), .A2(n6039), .B1(n6660), .B2(
        \registers[12][10] ), .ZN(n2605) );
  INV_X1 U2999 ( .A(n2604), .ZN(n3734) );
  AOI22_X1 U3000 ( .A1(datain[11]), .A2(n6039), .B1(n6662), .B2(
        \registers[12][11] ), .ZN(n2604) );
  INV_X1 U3001 ( .A(n2603), .ZN(n3735) );
  AOI22_X1 U3002 ( .A1(datain[12]), .A2(n6040), .B1(n6656), .B2(
        \registers[12][12] ), .ZN(n2603) );
  INV_X1 U3003 ( .A(n2602), .ZN(n3736) );
  AOI22_X1 U3004 ( .A1(datain[13]), .A2(n6040), .B1(n6657), .B2(
        \registers[12][13] ), .ZN(n2602) );
  INV_X1 U3005 ( .A(n2601), .ZN(n3737) );
  AOI22_X1 U3006 ( .A1(datain[14]), .A2(n6040), .B1(n6658), .B2(
        \registers[12][14] ), .ZN(n2601) );
  INV_X1 U3007 ( .A(n2600), .ZN(n3738) );
  AOI22_X1 U3008 ( .A1(datain[15]), .A2(n6040), .B1(n6657), .B2(
        \registers[12][15] ), .ZN(n2600) );
  INV_X1 U3009 ( .A(n2599), .ZN(n3739) );
  AOI22_X1 U3010 ( .A1(datain[16]), .A2(n6040), .B1(n6659), .B2(
        \registers[12][16] ), .ZN(n2599) );
  INV_X1 U3011 ( .A(n2598), .ZN(n3740) );
  AOI22_X1 U3012 ( .A1(datain[17]), .A2(n6040), .B1(n6659), .B2(
        \registers[12][17] ), .ZN(n2598) );
  INV_X1 U3013 ( .A(n2597), .ZN(n3741) );
  AOI22_X1 U3014 ( .A1(datain[18]), .A2(n6040), .B1(n6660), .B2(
        \registers[12][18] ), .ZN(n2597) );
  INV_X1 U3015 ( .A(n2596), .ZN(n3742) );
  AOI22_X1 U3016 ( .A1(datain[19]), .A2(n6040), .B1(n6659), .B2(
        \registers[12][19] ), .ZN(n2596) );
  INV_X1 U3017 ( .A(n2595), .ZN(n3743) );
  AOI22_X1 U3018 ( .A1(datain[20]), .A2(n6040), .B1(n6661), .B2(
        \registers[12][20] ), .ZN(n2595) );
  INV_X1 U3019 ( .A(n2594), .ZN(n3744) );
  AOI22_X1 U3020 ( .A1(datain[21]), .A2(n6040), .B1(n6662), .B2(
        \registers[12][21] ), .ZN(n2594) );
  INV_X1 U3021 ( .A(n2593), .ZN(n3745) );
  AOI22_X1 U3022 ( .A1(datain[22]), .A2(n6040), .B1(n6661), .B2(
        \registers[12][22] ), .ZN(n2593) );
  INV_X1 U3023 ( .A(n2592), .ZN(n3746) );
  AOI22_X1 U3024 ( .A1(datain[23]), .A2(n6040), .B1(n6661), .B2(
        \registers[12][23] ), .ZN(n2592) );
  INV_X1 U3025 ( .A(n2591), .ZN(n3747) );
  AOI22_X1 U3026 ( .A1(datain[24]), .A2(n6041), .B1(n6662), .B2(
        \registers[12][24] ), .ZN(n2591) );
  INV_X1 U3027 ( .A(n2590), .ZN(n3748) );
  AOI22_X1 U3028 ( .A1(datain[25]), .A2(n6041), .B1(n6662), .B2(
        \registers[12][25] ), .ZN(n2590) );
  INV_X1 U3029 ( .A(n2589), .ZN(n3749) );
  AOI22_X1 U3030 ( .A1(datain[26]), .A2(n6041), .B1(n6656), .B2(
        \registers[12][26] ), .ZN(n2589) );
  INV_X1 U3031 ( .A(n2588), .ZN(n3750) );
  AOI22_X1 U3032 ( .A1(datain[27]), .A2(n6041), .B1(n6656), .B2(
        \registers[12][27] ), .ZN(n2588) );
  INV_X1 U3033 ( .A(n2587), .ZN(n3751) );
  AOI22_X1 U3034 ( .A1(datain[28]), .A2(n6041), .B1(n6656), .B2(
        \registers[12][28] ), .ZN(n2587) );
  INV_X1 U3035 ( .A(n2586), .ZN(n3752) );
  AOI22_X1 U3036 ( .A1(datain[29]), .A2(n6041), .B1(n6662), .B2(
        \registers[12][29] ), .ZN(n2586) );
  INV_X1 U3037 ( .A(n2585), .ZN(n3753) );
  AOI22_X1 U3038 ( .A1(datain[30]), .A2(n6041), .B1(n6657), .B2(
        \registers[12][30] ), .ZN(n2585) );
  INV_X1 U3039 ( .A(n2582), .ZN(n3754) );
  AOI22_X1 U3040 ( .A1(datain[31]), .A2(n6041), .B1(n6660), .B2(
        \registers[12][31] ), .ZN(n2582) );
  INV_X1 U3041 ( .A(n1996), .ZN(n3883) );
  AOI22_X1 U3042 ( .A1(datain[0]), .A2(n6054), .B1(n6700), .B2(
        \registers[7][0] ), .ZN(n1996) );
  INV_X1 U3043 ( .A(n1995), .ZN(n3884) );
  AOI22_X1 U3044 ( .A1(datain[1]), .A2(n6054), .B1(n6701), .B2(
        \registers[7][1] ), .ZN(n1995) );
  INV_X1 U3045 ( .A(n1994), .ZN(n3885) );
  AOI22_X1 U3046 ( .A1(datain[2]), .A2(n6054), .B1(n6701), .B2(
        \registers[7][2] ), .ZN(n1994) );
  INV_X1 U3047 ( .A(n1993), .ZN(n3886) );
  AOI22_X1 U3048 ( .A1(datain[3]), .A2(n6054), .B1(n6700), .B2(
        \registers[7][3] ), .ZN(n1993) );
  INV_X1 U3049 ( .A(n1992), .ZN(n3887) );
  AOI22_X1 U3050 ( .A1(datain[4]), .A2(n6054), .B1(n6701), .B2(
        \registers[7][4] ), .ZN(n1992) );
  INV_X1 U3051 ( .A(n1991), .ZN(n3888) );
  AOI22_X1 U3052 ( .A1(datain[5]), .A2(n6054), .B1(n6702), .B2(
        \registers[7][5] ), .ZN(n1991) );
  INV_X1 U3053 ( .A(n1990), .ZN(n3889) );
  AOI22_X1 U3054 ( .A1(datain[6]), .A2(n6054), .B1(n6702), .B2(
        \registers[7][6] ), .ZN(n1990) );
  INV_X1 U3055 ( .A(n1989), .ZN(n3890) );
  AOI22_X1 U3056 ( .A1(datain[7]), .A2(n6054), .B1(n6703), .B2(
        \registers[7][7] ), .ZN(n1989) );
  INV_X1 U3057 ( .A(n1988), .ZN(n3891) );
  AOI22_X1 U3058 ( .A1(datain[8]), .A2(n6054), .B1(n6702), .B2(
        \registers[7][8] ), .ZN(n1988) );
  INV_X1 U3059 ( .A(n1987), .ZN(n3892) );
  AOI22_X1 U3060 ( .A1(datain[9]), .A2(n6054), .B1(n6703), .B2(
        \registers[7][9] ), .ZN(n1987) );
  INV_X1 U3061 ( .A(n1986), .ZN(n3893) );
  AOI22_X1 U3062 ( .A1(datain[10]), .A2(n6054), .B1(n6704), .B2(
        \registers[7][10] ), .ZN(n1986) );
  INV_X1 U3063 ( .A(n1985), .ZN(n3894) );
  AOI22_X1 U3064 ( .A1(datain[11]), .A2(n6054), .B1(n6705), .B2(
        \registers[7][11] ), .ZN(n1985) );
  INV_X1 U3065 ( .A(n1984), .ZN(n3895) );
  AOI22_X1 U3066 ( .A1(datain[12]), .A2(n6055), .B1(n6704), .B2(
        \registers[7][12] ), .ZN(n1984) );
  INV_X1 U3067 ( .A(n1983), .ZN(n3896) );
  AOI22_X1 U3068 ( .A1(datain[13]), .A2(n6055), .B1(n6705), .B2(
        \registers[7][13] ), .ZN(n1983) );
  INV_X1 U3069 ( .A(n1982), .ZN(n3897) );
  AOI22_X1 U3070 ( .A1(datain[14]), .A2(n6055), .B1(n6703), .B2(
        \registers[7][14] ), .ZN(n1982) );
  INV_X1 U3071 ( .A(n1981), .ZN(n3898) );
  AOI22_X1 U3072 ( .A1(datain[15]), .A2(n6055), .B1(n6700), .B2(
        \registers[7][15] ), .ZN(n1981) );
  INV_X1 U3073 ( .A(n1980), .ZN(n3899) );
  AOI22_X1 U3074 ( .A1(datain[16]), .A2(n6055), .B1(n6701), .B2(
        \registers[7][16] ), .ZN(n1980) );
  INV_X1 U3075 ( .A(n1979), .ZN(n3900) );
  AOI22_X1 U3076 ( .A1(datain[17]), .A2(n6055), .B1(n6702), .B2(
        \registers[7][17] ), .ZN(n1979) );
  INV_X1 U3077 ( .A(n1978), .ZN(n3901) );
  AOI22_X1 U3078 ( .A1(datain[18]), .A2(n6055), .B1(n6700), .B2(
        \registers[7][18] ), .ZN(n1978) );
  INV_X1 U3079 ( .A(n1977), .ZN(n3902) );
  AOI22_X1 U3080 ( .A1(datain[19]), .A2(n6055), .B1(n6701), .B2(
        \registers[7][19] ), .ZN(n1977) );
  INV_X1 U3081 ( .A(n1976), .ZN(n3903) );
  AOI22_X1 U3082 ( .A1(datain[20]), .A2(n6055), .B1(n6704), .B2(
        \registers[7][20] ), .ZN(n1976) );
  INV_X1 U3083 ( .A(n1975), .ZN(n3904) );
  AOI22_X1 U3084 ( .A1(datain[21]), .A2(n6055), .B1(n6703), .B2(
        \registers[7][21] ), .ZN(n1975) );
  INV_X1 U3085 ( .A(n1974), .ZN(n3905) );
  AOI22_X1 U3086 ( .A1(datain[22]), .A2(n6055), .B1(n6704), .B2(
        \registers[7][22] ), .ZN(n1974) );
  INV_X1 U3087 ( .A(n1973), .ZN(n3906) );
  AOI22_X1 U3088 ( .A1(datain[23]), .A2(n6055), .B1(n6705), .B2(
        \registers[7][23] ), .ZN(n1973) );
  INV_X1 U3089 ( .A(n1972), .ZN(n3907) );
  AOI22_X1 U3090 ( .A1(datain[24]), .A2(n6056), .B1(n6702), .B2(
        \registers[7][24] ), .ZN(n1972) );
  INV_X1 U3091 ( .A(n1971), .ZN(n3908) );
  AOI22_X1 U3092 ( .A1(datain[25]), .A2(n6056), .B1(n6703), .B2(
        \registers[7][25] ), .ZN(n1971) );
  INV_X1 U3093 ( .A(n1970), .ZN(n3909) );
  AOI22_X1 U3094 ( .A1(datain[26]), .A2(n6056), .B1(n6705), .B2(
        \registers[7][26] ), .ZN(n1970) );
  INV_X1 U3095 ( .A(n1969), .ZN(n3910) );
  AOI22_X1 U3096 ( .A1(datain[27]), .A2(n6056), .B1(n6700), .B2(
        \registers[7][27] ), .ZN(n1969) );
  INV_X1 U3097 ( .A(n1968), .ZN(n3911) );
  AOI22_X1 U3098 ( .A1(datain[28]), .A2(n6056), .B1(n6701), .B2(
        \registers[7][28] ), .ZN(n1968) );
  INV_X1 U3099 ( .A(n1967), .ZN(n3912) );
  AOI22_X1 U3100 ( .A1(datain[29]), .A2(n6056), .B1(n6702), .B2(
        \registers[7][29] ), .ZN(n1967) );
  INV_X1 U3101 ( .A(n1966), .ZN(n3913) );
  AOI22_X1 U3102 ( .A1(datain[30]), .A2(n6056), .B1(n6704), .B2(
        \registers[7][30] ), .ZN(n1966) );
  INV_X1 U3103 ( .A(n1963), .ZN(n3914) );
  AOI22_X1 U3104 ( .A1(datain[31]), .A2(n6056), .B1(n6705), .B2(
        \registers[7][31] ), .ZN(n1963) );
  INV_X1 U3105 ( .A(n1962), .ZN(n3915) );
  AOI22_X1 U3106 ( .A1(datain[0]), .A2(n6057), .B1(n6707), .B2(
        \registers[6][0] ), .ZN(n1962) );
  INV_X1 U3107 ( .A(n1961), .ZN(n3916) );
  AOI22_X1 U3108 ( .A1(datain[1]), .A2(n6057), .B1(n6708), .B2(
        \registers[6][1] ), .ZN(n1961) );
  INV_X1 U3109 ( .A(n1960), .ZN(n3917) );
  AOI22_X1 U3110 ( .A1(datain[2]), .A2(n6057), .B1(n6708), .B2(
        \registers[6][2] ), .ZN(n1960) );
  INV_X1 U3111 ( .A(n1959), .ZN(n3918) );
  AOI22_X1 U3112 ( .A1(datain[3]), .A2(n6057), .B1(n6707), .B2(
        \registers[6][3] ), .ZN(n1959) );
  INV_X1 U3113 ( .A(n1958), .ZN(n3919) );
  AOI22_X1 U3114 ( .A1(datain[4]), .A2(n6057), .B1(n6708), .B2(
        \registers[6][4] ), .ZN(n1958) );
  INV_X1 U3115 ( .A(n1957), .ZN(n3920) );
  AOI22_X1 U3116 ( .A1(datain[5]), .A2(n6057), .B1(n6709), .B2(
        \registers[6][5] ), .ZN(n1957) );
  INV_X1 U3117 ( .A(n1956), .ZN(n3921) );
  AOI22_X1 U3118 ( .A1(datain[6]), .A2(n6057), .B1(n6709), .B2(
        \registers[6][6] ), .ZN(n1956) );
  INV_X1 U3119 ( .A(n1955), .ZN(n3922) );
  AOI22_X1 U3120 ( .A1(datain[7]), .A2(n6057), .B1(n6710), .B2(
        \registers[6][7] ), .ZN(n1955) );
  INV_X1 U3121 ( .A(n1954), .ZN(n3923) );
  AOI22_X1 U3122 ( .A1(datain[8]), .A2(n6057), .B1(n6709), .B2(
        \registers[6][8] ), .ZN(n1954) );
  INV_X1 U3123 ( .A(n1953), .ZN(n3924) );
  AOI22_X1 U3124 ( .A1(datain[9]), .A2(n6057), .B1(n6710), .B2(
        \registers[6][9] ), .ZN(n1953) );
  INV_X1 U3125 ( .A(n1952), .ZN(n3925) );
  AOI22_X1 U3126 ( .A1(datain[10]), .A2(n6057), .B1(n6711), .B2(
        \registers[6][10] ), .ZN(n1952) );
  INV_X1 U3127 ( .A(n1951), .ZN(n3926) );
  AOI22_X1 U3128 ( .A1(datain[11]), .A2(n6057), .B1(n6712), .B2(
        \registers[6][11] ), .ZN(n1951) );
  INV_X1 U3129 ( .A(n1950), .ZN(n3927) );
  AOI22_X1 U3130 ( .A1(datain[12]), .A2(n6058), .B1(n6711), .B2(
        \registers[6][12] ), .ZN(n1950) );
  INV_X1 U3131 ( .A(n1949), .ZN(n3928) );
  AOI22_X1 U3132 ( .A1(datain[13]), .A2(n6058), .B1(n6712), .B2(
        \registers[6][13] ), .ZN(n1949) );
  INV_X1 U3133 ( .A(n1948), .ZN(n3929) );
  AOI22_X1 U3134 ( .A1(datain[14]), .A2(n6058), .B1(n6710), .B2(
        \registers[6][14] ), .ZN(n1948) );
  INV_X1 U3135 ( .A(n1947), .ZN(n3930) );
  AOI22_X1 U3136 ( .A1(datain[15]), .A2(n6058), .B1(n6707), .B2(
        \registers[6][15] ), .ZN(n1947) );
  INV_X1 U3137 ( .A(n1946), .ZN(n3931) );
  AOI22_X1 U3138 ( .A1(datain[16]), .A2(n6058), .B1(n6708), .B2(
        \registers[6][16] ), .ZN(n1946) );
  INV_X1 U3139 ( .A(n1945), .ZN(n3932) );
  AOI22_X1 U3140 ( .A1(datain[17]), .A2(n6058), .B1(n6709), .B2(
        \registers[6][17] ), .ZN(n1945) );
  INV_X1 U3141 ( .A(n1944), .ZN(n3933) );
  AOI22_X1 U3142 ( .A1(datain[18]), .A2(n6058), .B1(n6707), .B2(
        \registers[6][18] ), .ZN(n1944) );
  INV_X1 U3143 ( .A(n1943), .ZN(n3934) );
  AOI22_X1 U3144 ( .A1(datain[19]), .A2(n6058), .B1(n6708), .B2(
        \registers[6][19] ), .ZN(n1943) );
  INV_X1 U3145 ( .A(n1942), .ZN(n3935) );
  AOI22_X1 U3146 ( .A1(datain[20]), .A2(n6058), .B1(n6711), .B2(
        \registers[6][20] ), .ZN(n1942) );
  INV_X1 U3147 ( .A(n1941), .ZN(n3936) );
  AOI22_X1 U3148 ( .A1(datain[21]), .A2(n6058), .B1(n6710), .B2(
        \registers[6][21] ), .ZN(n1941) );
  INV_X1 U3149 ( .A(n1940), .ZN(n3937) );
  AOI22_X1 U3150 ( .A1(datain[22]), .A2(n6058), .B1(n6711), .B2(
        \registers[6][22] ), .ZN(n1940) );
  INV_X1 U3151 ( .A(n1939), .ZN(n3938) );
  AOI22_X1 U3152 ( .A1(datain[23]), .A2(n6058), .B1(n6712), .B2(
        \registers[6][23] ), .ZN(n1939) );
  INV_X1 U3153 ( .A(n1938), .ZN(n3939) );
  AOI22_X1 U3154 ( .A1(datain[24]), .A2(n6059), .B1(n6709), .B2(
        \registers[6][24] ), .ZN(n1938) );
  INV_X1 U3155 ( .A(n1937), .ZN(n3940) );
  AOI22_X1 U3156 ( .A1(datain[25]), .A2(n6059), .B1(n6710), .B2(
        \registers[6][25] ), .ZN(n1937) );
  INV_X1 U3157 ( .A(n1936), .ZN(n3941) );
  AOI22_X1 U3158 ( .A1(datain[26]), .A2(n6059), .B1(n6712), .B2(
        \registers[6][26] ), .ZN(n1936) );
  INV_X1 U3159 ( .A(n1935), .ZN(n3942) );
  AOI22_X1 U3160 ( .A1(datain[27]), .A2(n6059), .B1(n6707), .B2(
        \registers[6][27] ), .ZN(n1935) );
  INV_X1 U3161 ( .A(n1934), .ZN(n3943) );
  AOI22_X1 U3162 ( .A1(datain[28]), .A2(n6059), .B1(n6708), .B2(
        \registers[6][28] ), .ZN(n1934) );
  INV_X1 U3163 ( .A(n1933), .ZN(n3944) );
  AOI22_X1 U3164 ( .A1(datain[29]), .A2(n6059), .B1(n6709), .B2(
        \registers[6][29] ), .ZN(n1933) );
  INV_X1 U3165 ( .A(n1932), .ZN(n3945) );
  AOI22_X1 U3166 ( .A1(datain[30]), .A2(n6059), .B1(n6711), .B2(
        \registers[6][30] ), .ZN(n1932) );
  INV_X1 U3167 ( .A(n1929), .ZN(n3946) );
  AOI22_X1 U3168 ( .A1(datain[31]), .A2(n6059), .B1(n6712), .B2(
        \registers[6][31] ), .ZN(n1929) );
  INV_X1 U3169 ( .A(n1928), .ZN(n3947) );
  AOI22_X1 U3170 ( .A1(datain[0]), .A2(n6060), .B1(n6715), .B2(
        \registers[5][0] ), .ZN(n1928) );
  INV_X1 U3171 ( .A(n1927), .ZN(n3948) );
  AOI22_X1 U3172 ( .A1(datain[1]), .A2(n6060), .B1(n6716), .B2(
        \registers[5][1] ), .ZN(n1927) );
  INV_X1 U3173 ( .A(n1926), .ZN(n3949) );
  AOI22_X1 U3174 ( .A1(datain[2]), .A2(n6060), .B1(n6717), .B2(
        \registers[5][2] ), .ZN(n1926) );
  INV_X1 U3175 ( .A(n1925), .ZN(n3950) );
  AOI22_X1 U3176 ( .A1(datain[3]), .A2(n6060), .B1(n6720), .B2(
        \registers[5][3] ), .ZN(n1925) );
  INV_X1 U3177 ( .A(n1924), .ZN(n3951) );
  AOI22_X1 U3178 ( .A1(datain[4]), .A2(n6060), .B1(n6716), .B2(
        \registers[5][4] ), .ZN(n1924) );
  INV_X1 U3179 ( .A(n1923), .ZN(n3952) );
  AOI22_X1 U3180 ( .A1(datain[5]), .A2(n6060), .B1(n6717), .B2(
        \registers[5][5] ), .ZN(n1923) );
  INV_X1 U3181 ( .A(n1922), .ZN(n3953) );
  AOI22_X1 U3182 ( .A1(datain[6]), .A2(n6060), .B1(n6717), .B2(
        \registers[5][6] ), .ZN(n1922) );
  INV_X1 U3183 ( .A(n1921), .ZN(n3954) );
  AOI22_X1 U3184 ( .A1(datain[7]), .A2(n6060), .B1(n6718), .B2(
        \registers[5][7] ), .ZN(n1921) );
  INV_X1 U3185 ( .A(n1920), .ZN(n3955) );
  AOI22_X1 U3186 ( .A1(datain[8]), .A2(n6060), .B1(n6718), .B2(
        \registers[5][8] ), .ZN(n1920) );
  INV_X1 U3187 ( .A(n1919), .ZN(n3956) );
  AOI22_X1 U3188 ( .A1(datain[9]), .A2(n6060), .B1(n6719), .B2(
        \registers[5][9] ), .ZN(n1919) );
  INV_X1 U3189 ( .A(n1918), .ZN(n3957) );
  AOI22_X1 U3190 ( .A1(datain[10]), .A2(n6060), .B1(n6719), .B2(
        \registers[5][10] ), .ZN(n1918) );
  INV_X1 U3191 ( .A(n1917), .ZN(n3958) );
  AOI22_X1 U3192 ( .A1(datain[11]), .A2(n6060), .B1(n6721), .B2(
        \registers[5][11] ), .ZN(n1917) );
  INV_X1 U3193 ( .A(n1916), .ZN(n3959) );
  AOI22_X1 U3194 ( .A1(datain[12]), .A2(n6061), .B1(n6715), .B2(
        \registers[5][12] ), .ZN(n1916) );
  INV_X1 U3195 ( .A(n1915), .ZN(n3960) );
  AOI22_X1 U3196 ( .A1(datain[13]), .A2(n6061), .B1(n6716), .B2(
        \registers[5][13] ), .ZN(n1915) );
  INV_X1 U3197 ( .A(n1914), .ZN(n3961) );
  AOI22_X1 U3198 ( .A1(datain[14]), .A2(n6061), .B1(n6717), .B2(
        \registers[5][14] ), .ZN(n1914) );
  INV_X1 U3199 ( .A(n1913), .ZN(n3962) );
  AOI22_X1 U3200 ( .A1(datain[15]), .A2(n6061), .B1(n6716), .B2(
        \registers[5][15] ), .ZN(n1913) );
  INV_X1 U3201 ( .A(n1912), .ZN(n3963) );
  AOI22_X1 U3202 ( .A1(datain[16]), .A2(n6061), .B1(n6718), .B2(
        \registers[5][16] ), .ZN(n1912) );
  INV_X1 U3203 ( .A(n1911), .ZN(n3964) );
  AOI22_X1 U3204 ( .A1(datain[17]), .A2(n6061), .B1(n6718), .B2(
        \registers[5][17] ), .ZN(n1911) );
  INV_X1 U3205 ( .A(n1910), .ZN(n3965) );
  AOI22_X1 U3206 ( .A1(datain[18]), .A2(n6061), .B1(n6719), .B2(
        \registers[5][18] ), .ZN(n1910) );
  INV_X1 U3207 ( .A(n1909), .ZN(n3966) );
  AOI22_X1 U3208 ( .A1(datain[19]), .A2(n6061), .B1(n6718), .B2(
        \registers[5][19] ), .ZN(n1909) );
  INV_X1 U3209 ( .A(n1908), .ZN(n3967) );
  AOI22_X1 U3210 ( .A1(datain[20]), .A2(n6061), .B1(n6720), .B2(
        \registers[5][20] ), .ZN(n1908) );
  INV_X1 U3211 ( .A(n1907), .ZN(n3968) );
  AOI22_X1 U3212 ( .A1(datain[21]), .A2(n6061), .B1(n6721), .B2(
        \registers[5][21] ), .ZN(n1907) );
  INV_X1 U3213 ( .A(n1906), .ZN(n3969) );
  AOI22_X1 U3214 ( .A1(datain[22]), .A2(n6061), .B1(n6720), .B2(
        \registers[5][22] ), .ZN(n1906) );
  INV_X1 U3215 ( .A(n1905), .ZN(n3970) );
  AOI22_X1 U3216 ( .A1(datain[23]), .A2(n6061), .B1(n6720), .B2(
        \registers[5][23] ), .ZN(n1905) );
  INV_X1 U3217 ( .A(n1904), .ZN(n3971) );
  AOI22_X1 U3218 ( .A1(datain[24]), .A2(n6062), .B1(n6721), .B2(
        \registers[5][24] ), .ZN(n1904) );
  INV_X1 U3219 ( .A(n1903), .ZN(n3972) );
  AOI22_X1 U3220 ( .A1(datain[25]), .A2(n6062), .B1(n6721), .B2(
        \registers[5][25] ), .ZN(n1903) );
  INV_X1 U3221 ( .A(n1902), .ZN(n3973) );
  AOI22_X1 U3222 ( .A1(datain[26]), .A2(n6062), .B1(n6715), .B2(
        \registers[5][26] ), .ZN(n1902) );
  INV_X1 U3223 ( .A(n1901), .ZN(n3974) );
  AOI22_X1 U3224 ( .A1(datain[27]), .A2(n6062), .B1(n6715), .B2(
        \registers[5][27] ), .ZN(n1901) );
  INV_X1 U3225 ( .A(n1900), .ZN(n3975) );
  AOI22_X1 U3226 ( .A1(datain[28]), .A2(n6062), .B1(n6715), .B2(
        \registers[5][28] ), .ZN(n1900) );
  INV_X1 U3227 ( .A(n1899), .ZN(n3976) );
  AOI22_X1 U3228 ( .A1(datain[29]), .A2(n6062), .B1(n6721), .B2(
        \registers[5][29] ), .ZN(n1899) );
  INV_X1 U3229 ( .A(n1898), .ZN(n3977) );
  AOI22_X1 U3230 ( .A1(datain[30]), .A2(n6062), .B1(n6716), .B2(
        \registers[5][30] ), .ZN(n1898) );
  INV_X1 U3231 ( .A(n1895), .ZN(n3978) );
  AOI22_X1 U3232 ( .A1(datain[31]), .A2(n6062), .B1(n6719), .B2(
        \registers[5][31] ), .ZN(n1895) );
  INV_X1 U3233 ( .A(n1893), .ZN(n3979) );
  AOI22_X1 U3234 ( .A1(datain[0]), .A2(n6063), .B1(n6724), .B2(
        \registers[4][0] ), .ZN(n1893) );
  INV_X1 U3235 ( .A(n1892), .ZN(n3980) );
  AOI22_X1 U3236 ( .A1(datain[1]), .A2(n6063), .B1(n6725), .B2(
        \registers[4][1] ), .ZN(n1892) );
  INV_X1 U3237 ( .A(n1891), .ZN(n3981) );
  AOI22_X1 U3238 ( .A1(datain[2]), .A2(n6063), .B1(n6726), .B2(
        \registers[4][2] ), .ZN(n1891) );
  INV_X1 U3239 ( .A(n1890), .ZN(n3982) );
  AOI22_X1 U3240 ( .A1(datain[3]), .A2(n6063), .B1(n6729), .B2(
        \registers[4][3] ), .ZN(n1890) );
  INV_X1 U3241 ( .A(n1889), .ZN(n3983) );
  AOI22_X1 U3242 ( .A1(datain[4]), .A2(n6063), .B1(n6725), .B2(
        \registers[4][4] ), .ZN(n1889) );
  INV_X1 U3243 ( .A(n1888), .ZN(n3984) );
  AOI22_X1 U3244 ( .A1(datain[5]), .A2(n6063), .B1(n6726), .B2(
        \registers[4][5] ), .ZN(n1888) );
  INV_X1 U3245 ( .A(n1887), .ZN(n3985) );
  AOI22_X1 U3246 ( .A1(datain[6]), .A2(n6063), .B1(n6726), .B2(
        \registers[4][6] ), .ZN(n1887) );
  INV_X1 U3247 ( .A(n1886), .ZN(n3986) );
  AOI22_X1 U3248 ( .A1(datain[7]), .A2(n6063), .B1(n6727), .B2(
        \registers[4][7] ), .ZN(n1886) );
  INV_X1 U3249 ( .A(n1885), .ZN(n3987) );
  AOI22_X1 U3250 ( .A1(datain[8]), .A2(n6063), .B1(n6727), .B2(
        \registers[4][8] ), .ZN(n1885) );
  INV_X1 U3251 ( .A(n1884), .ZN(n3988) );
  AOI22_X1 U3252 ( .A1(datain[9]), .A2(n6063), .B1(n6728), .B2(
        \registers[4][9] ), .ZN(n1884) );
  INV_X1 U3253 ( .A(n1883), .ZN(n3989) );
  AOI22_X1 U3254 ( .A1(datain[10]), .A2(n6063), .B1(n6728), .B2(
        \registers[4][10] ), .ZN(n1883) );
  INV_X1 U3255 ( .A(n1882), .ZN(n3990) );
  AOI22_X1 U3256 ( .A1(datain[11]), .A2(n6063), .B1(n6730), .B2(
        \registers[4][11] ), .ZN(n1882) );
  INV_X1 U3257 ( .A(n1881), .ZN(n3991) );
  AOI22_X1 U3258 ( .A1(datain[12]), .A2(n6064), .B1(n6724), .B2(
        \registers[4][12] ), .ZN(n1881) );
  INV_X1 U3259 ( .A(n1880), .ZN(n3992) );
  AOI22_X1 U3260 ( .A1(datain[13]), .A2(n6064), .B1(n6725), .B2(
        \registers[4][13] ), .ZN(n1880) );
  INV_X1 U3261 ( .A(n1879), .ZN(n3993) );
  AOI22_X1 U3262 ( .A1(datain[14]), .A2(n6064), .B1(n6726), .B2(
        \registers[4][14] ), .ZN(n1879) );
  INV_X1 U3263 ( .A(n1878), .ZN(n3994) );
  AOI22_X1 U3264 ( .A1(datain[15]), .A2(n6064), .B1(n6725), .B2(
        \registers[4][15] ), .ZN(n1878) );
  INV_X1 U3265 ( .A(n1877), .ZN(n3995) );
  AOI22_X1 U3266 ( .A1(datain[16]), .A2(n6064), .B1(n6727), .B2(
        \registers[4][16] ), .ZN(n1877) );
  INV_X1 U3267 ( .A(n1876), .ZN(n3996) );
  AOI22_X1 U3268 ( .A1(datain[17]), .A2(n6064), .B1(n6727), .B2(
        \registers[4][17] ), .ZN(n1876) );
  INV_X1 U3269 ( .A(n1875), .ZN(n3997) );
  AOI22_X1 U3270 ( .A1(datain[18]), .A2(n6064), .B1(n6728), .B2(
        \registers[4][18] ), .ZN(n1875) );
  INV_X1 U3271 ( .A(n1874), .ZN(n3998) );
  AOI22_X1 U3272 ( .A1(datain[19]), .A2(n6064), .B1(n6727), .B2(
        \registers[4][19] ), .ZN(n1874) );
  INV_X1 U3273 ( .A(n1873), .ZN(n3999) );
  AOI22_X1 U3274 ( .A1(datain[20]), .A2(n6064), .B1(n6729), .B2(
        \registers[4][20] ), .ZN(n1873) );
  INV_X1 U3275 ( .A(n1872), .ZN(n4000) );
  AOI22_X1 U3276 ( .A1(datain[21]), .A2(n6064), .B1(n6730), .B2(
        \registers[4][21] ), .ZN(n1872) );
  INV_X1 U3277 ( .A(n1871), .ZN(n4001) );
  AOI22_X1 U3278 ( .A1(datain[22]), .A2(n6064), .B1(n6729), .B2(
        \registers[4][22] ), .ZN(n1871) );
  INV_X1 U3279 ( .A(n1870), .ZN(n4002) );
  AOI22_X1 U3280 ( .A1(datain[23]), .A2(n6064), .B1(n6729), .B2(
        \registers[4][23] ), .ZN(n1870) );
  INV_X1 U3281 ( .A(n1869), .ZN(n4003) );
  AOI22_X1 U3282 ( .A1(datain[24]), .A2(n6065), .B1(n6730), .B2(
        \registers[4][24] ), .ZN(n1869) );
  INV_X1 U3283 ( .A(n1868), .ZN(n4004) );
  AOI22_X1 U3284 ( .A1(datain[25]), .A2(n6065), .B1(n6730), .B2(
        \registers[4][25] ), .ZN(n1868) );
  INV_X1 U3285 ( .A(n1867), .ZN(n4005) );
  AOI22_X1 U3286 ( .A1(datain[26]), .A2(n6065), .B1(n6724), .B2(
        \registers[4][26] ), .ZN(n1867) );
  INV_X1 U3287 ( .A(n1866), .ZN(n4006) );
  AOI22_X1 U3288 ( .A1(datain[27]), .A2(n6065), .B1(n6724), .B2(
        \registers[4][27] ), .ZN(n1866) );
  INV_X1 U3289 ( .A(n1865), .ZN(n4007) );
  AOI22_X1 U3290 ( .A1(datain[28]), .A2(n6065), .B1(n6724), .B2(
        \registers[4][28] ), .ZN(n1865) );
  INV_X1 U3291 ( .A(n1864), .ZN(n4008) );
  AOI22_X1 U3292 ( .A1(datain[29]), .A2(n6065), .B1(n6730), .B2(
        \registers[4][29] ), .ZN(n1864) );
  INV_X1 U3293 ( .A(n1863), .ZN(n4009) );
  AOI22_X1 U3294 ( .A1(datain[30]), .A2(n6065), .B1(n6725), .B2(
        \registers[4][30] ), .ZN(n1863) );
  INV_X1 U3295 ( .A(n1860), .ZN(n4010) );
  AOI22_X1 U3296 ( .A1(datain[31]), .A2(n6065), .B1(n6728), .B2(
        \registers[4][31] ), .ZN(n1860) );
  INV_X1 U3297 ( .A(enable), .ZN(n2719) );
  INV_X1 U3298 ( .A(n5140), .ZN(n6076) );
  INV_X1 U3299 ( .A(n6076), .ZN(n6077) );
  INV_X1 U3300 ( .A(n6076), .ZN(n6078) );
  INV_X1 U3301 ( .A(n6076), .ZN(n6079) );
  INV_X1 U3302 ( .A(n6076), .ZN(n6080) );
  INV_X1 U3303 ( .A(n6076), .ZN(n6081) );
  INV_X1 U3304 ( .A(n6076), .ZN(n6082) );
  INV_X1 U3305 ( .A(n6076), .ZN(n6083) );
  INV_X1 U3306 ( .A(n5141), .ZN(n6084) );
  INV_X1 U3307 ( .A(n6084), .ZN(n6085) );
  INV_X1 U3308 ( .A(n6084), .ZN(n6086) );
  INV_X1 U3309 ( .A(n6084), .ZN(n6087) );
  INV_X1 U3310 ( .A(n6084), .ZN(n6088) );
  INV_X1 U3311 ( .A(n6084), .ZN(n6089) );
  INV_X1 U3312 ( .A(n6084), .ZN(n6090) );
  INV_X1 U3313 ( .A(n6084), .ZN(n6091) );
  INV_X1 U3314 ( .A(n6092), .ZN(n6093) );
  INV_X1 U3315 ( .A(n6092), .ZN(n6094) );
  INV_X1 U3316 ( .A(n6092), .ZN(n6095) );
  INV_X1 U3317 ( .A(n6092), .ZN(n6096) );
  INV_X1 U3318 ( .A(n6092), .ZN(n6097) );
  INV_X1 U3319 ( .A(n6092), .ZN(n6098) );
  INV_X1 U3320 ( .A(n6092), .ZN(n6099) );
  INV_X1 U3321 ( .A(n6100), .ZN(n6101) );
  INV_X1 U3322 ( .A(n6100), .ZN(n6102) );
  INV_X1 U3323 ( .A(n6100), .ZN(n6103) );
  INV_X1 U3324 ( .A(n6100), .ZN(n6104) );
  INV_X1 U3325 ( .A(n6100), .ZN(n6105) );
  INV_X1 U3326 ( .A(n6100), .ZN(n6106) );
  INV_X1 U3327 ( .A(n6100), .ZN(n6107) );
  INV_X1 U3328 ( .A(n5135), .ZN(n6108) );
  INV_X1 U3329 ( .A(n6108), .ZN(n6109) );
  INV_X1 U3330 ( .A(n6108), .ZN(n6110) );
  INV_X1 U3331 ( .A(n6108), .ZN(n6111) );
  INV_X1 U3332 ( .A(n6108), .ZN(n6112) );
  INV_X1 U3333 ( .A(n6108), .ZN(n6113) );
  INV_X1 U3334 ( .A(n6108), .ZN(n6114) );
  INV_X1 U3335 ( .A(n6108), .ZN(n6115) );
  INV_X1 U3336 ( .A(n6119), .ZN(n6120) );
  INV_X1 U3337 ( .A(n6119), .ZN(n6121) );
  INV_X1 U3338 ( .A(n6119), .ZN(n6122) );
  INV_X1 U3339 ( .A(n6119), .ZN(n6123) );
  INV_X1 U3340 ( .A(n6119), .ZN(n6124) );
  INV_X1 U3341 ( .A(n6119), .ZN(n6125) );
  INV_X1 U3342 ( .A(n6119), .ZN(n6126) );
  INV_X1 U3343 ( .A(n6127), .ZN(n6128) );
  INV_X1 U3344 ( .A(n6127), .ZN(n6129) );
  INV_X1 U3345 ( .A(n6127), .ZN(n6130) );
  INV_X1 U3346 ( .A(n6127), .ZN(n6131) );
  INV_X1 U3347 ( .A(n6127), .ZN(n6132) );
  INV_X1 U3348 ( .A(n6127), .ZN(n6133) );
  INV_X1 U3349 ( .A(n6127), .ZN(n6134) );
  INV_X1 U3350 ( .A(n5130), .ZN(n6135) );
  INV_X1 U3351 ( .A(n6135), .ZN(n6136) );
  INV_X1 U3352 ( .A(n6135), .ZN(n6137) );
  INV_X1 U3353 ( .A(n6135), .ZN(n6138) );
  INV_X1 U3354 ( .A(n6135), .ZN(n6139) );
  INV_X1 U3355 ( .A(n6135), .ZN(n6140) );
  INV_X1 U3356 ( .A(n6135), .ZN(n6141) );
  INV_X1 U3357 ( .A(n6135), .ZN(n6142) );
  INV_X1 U3358 ( .A(n6146), .ZN(n6147) );
  INV_X1 U3359 ( .A(n6146), .ZN(n6148) );
  INV_X1 U3360 ( .A(n6146), .ZN(n6149) );
  INV_X1 U3361 ( .A(n6146), .ZN(n6150) );
  INV_X1 U3362 ( .A(n6146), .ZN(n6151) );
  INV_X1 U3363 ( .A(n6146), .ZN(n6152) );
  INV_X1 U3364 ( .A(n6146), .ZN(n6153) );
  INV_X1 U3365 ( .A(n6154), .ZN(n6155) );
  INV_X1 U3366 ( .A(n6154), .ZN(n6156) );
  INV_X1 U3367 ( .A(n6154), .ZN(n6157) );
  INV_X1 U3368 ( .A(n6154), .ZN(n6158) );
  INV_X1 U3369 ( .A(n6154), .ZN(n6159) );
  INV_X1 U3370 ( .A(n6154), .ZN(n6160) );
  INV_X1 U3371 ( .A(n6154), .ZN(n6161) );
  INV_X1 U3372 ( .A(n5125), .ZN(n6162) );
  INV_X1 U3373 ( .A(n6162), .ZN(n6163) );
  INV_X1 U3374 ( .A(n6162), .ZN(n6164) );
  INV_X1 U3375 ( .A(n6162), .ZN(n6165) );
  INV_X1 U3376 ( .A(n6162), .ZN(n6166) );
  INV_X1 U3377 ( .A(n6162), .ZN(n6167) );
  INV_X1 U3378 ( .A(n6162), .ZN(n6168) );
  INV_X1 U3379 ( .A(n6162), .ZN(n6169) );
  INV_X1 U3380 ( .A(n6186), .ZN(n6187) );
  INV_X1 U3381 ( .A(n6186), .ZN(n6188) );
  INV_X1 U3382 ( .A(n6186), .ZN(n6189) );
  INV_X1 U3383 ( .A(n6186), .ZN(n6190) );
  INV_X1 U3384 ( .A(n6186), .ZN(n6191) );
  INV_X1 U3385 ( .A(n6186), .ZN(n6192) );
  INV_X1 U3386 ( .A(n6186), .ZN(n6193) );
  INV_X1 U3387 ( .A(n6194), .ZN(n6195) );
  INV_X1 U3388 ( .A(n6194), .ZN(n6196) );
  INV_X1 U3389 ( .A(n6194), .ZN(n6197) );
  INV_X1 U3390 ( .A(n6194), .ZN(n6198) );
  INV_X1 U3391 ( .A(n6194), .ZN(n6199) );
  INV_X1 U3392 ( .A(n6194), .ZN(n6200) );
  INV_X1 U3393 ( .A(n6194), .ZN(n6201) );
  INV_X1 U3394 ( .A(n5111), .ZN(n6202) );
  INV_X1 U3395 ( .A(n6202), .ZN(n6203) );
  INV_X1 U3396 ( .A(n6202), .ZN(n6204) );
  INV_X1 U3397 ( .A(n6202), .ZN(n6205) );
  INV_X1 U3398 ( .A(n6202), .ZN(n6206) );
  INV_X1 U3399 ( .A(n6202), .ZN(n6207) );
  INV_X1 U3400 ( .A(n6202), .ZN(n6208) );
  INV_X1 U3401 ( .A(n6202), .ZN(n6209) );
  INV_X1 U3402 ( .A(n5112), .ZN(n6210) );
  INV_X1 U3403 ( .A(n6210), .ZN(n6211) );
  INV_X1 U3404 ( .A(n6210), .ZN(n6212) );
  INV_X1 U3405 ( .A(n6210), .ZN(n6213) );
  INV_X1 U3406 ( .A(n6210), .ZN(n6214) );
  INV_X1 U3407 ( .A(n6210), .ZN(n6215) );
  INV_X1 U3408 ( .A(n6210), .ZN(n6216) );
  INV_X1 U3409 ( .A(n6210), .ZN(n6217) );
  INV_X1 U3410 ( .A(n6218), .ZN(n6219) );
  INV_X1 U3411 ( .A(n6218), .ZN(n6220) );
  INV_X1 U3412 ( .A(n6218), .ZN(n6221) );
  INV_X1 U3413 ( .A(n6218), .ZN(n6222) );
  INV_X1 U3414 ( .A(n6218), .ZN(n6223) );
  INV_X1 U3415 ( .A(n6218), .ZN(n6224) );
  INV_X1 U3416 ( .A(n6218), .ZN(n6225) );
  INV_X1 U3417 ( .A(n6226), .ZN(n6227) );
  INV_X1 U3418 ( .A(n6226), .ZN(n6228) );
  INV_X1 U3419 ( .A(n6226), .ZN(n6229) );
  INV_X1 U3420 ( .A(n6226), .ZN(n6230) );
  INV_X1 U3421 ( .A(n6226), .ZN(n6231) );
  INV_X1 U3422 ( .A(n6226), .ZN(n6232) );
  INV_X1 U3423 ( .A(n6226), .ZN(n6233) );
  INV_X1 U3424 ( .A(n5106), .ZN(n6234) );
  INV_X1 U3425 ( .A(n6234), .ZN(n6235) );
  INV_X1 U3426 ( .A(n6234), .ZN(n6236) );
  INV_X1 U3427 ( .A(n6234), .ZN(n6237) );
  INV_X1 U3428 ( .A(n6234), .ZN(n6238) );
  INV_X1 U3429 ( .A(n6234), .ZN(n6239) );
  INV_X1 U3430 ( .A(n6234), .ZN(n6240) );
  INV_X1 U3431 ( .A(n6234), .ZN(n6241) );
  INV_X1 U3432 ( .A(n6245), .ZN(n6246) );
  INV_X1 U3433 ( .A(n6245), .ZN(n6247) );
  INV_X1 U3434 ( .A(n6245), .ZN(n6248) );
  INV_X1 U3435 ( .A(n6245), .ZN(n6249) );
  INV_X1 U3436 ( .A(n6245), .ZN(n6250) );
  INV_X1 U3437 ( .A(n6245), .ZN(n6251) );
  INV_X1 U3438 ( .A(n6245), .ZN(n6252) );
  INV_X1 U3439 ( .A(n6253), .ZN(n6254) );
  INV_X1 U3440 ( .A(n6253), .ZN(n6255) );
  INV_X1 U3441 ( .A(n6253), .ZN(n6256) );
  INV_X1 U3442 ( .A(n6253), .ZN(n6257) );
  INV_X1 U3443 ( .A(n6253), .ZN(n6258) );
  INV_X1 U3444 ( .A(n6253), .ZN(n6259) );
  INV_X1 U3445 ( .A(n6253), .ZN(n6260) );
  INV_X1 U3446 ( .A(n4441), .ZN(n6281) );
  INV_X1 U3447 ( .A(n6281), .ZN(n6282) );
  INV_X1 U3448 ( .A(n6281), .ZN(n6283) );
  INV_X1 U3449 ( .A(n6281), .ZN(n6284) );
  INV_X1 U3450 ( .A(n6281), .ZN(n6285) );
  INV_X1 U3451 ( .A(n6281), .ZN(n6286) );
  INV_X1 U3452 ( .A(n6281), .ZN(n6287) );
  INV_X1 U3453 ( .A(n6281), .ZN(n6288) );
  INV_X1 U3454 ( .A(n6292), .ZN(n6293) );
  INV_X1 U3455 ( .A(n6292), .ZN(n6294) );
  INV_X1 U3456 ( .A(n6292), .ZN(n6295) );
  INV_X1 U3457 ( .A(n6292), .ZN(n6296) );
  INV_X1 U3458 ( .A(n6292), .ZN(n6297) );
  INV_X1 U3459 ( .A(n6292), .ZN(n6298) );
  INV_X1 U3460 ( .A(n6292), .ZN(n6299) );
  INV_X1 U3461 ( .A(n6300), .ZN(n6301) );
  INV_X1 U3462 ( .A(n6300), .ZN(n6302) );
  INV_X1 U3463 ( .A(n6300), .ZN(n6303) );
  INV_X1 U3464 ( .A(n6300), .ZN(n6304) );
  INV_X1 U3465 ( .A(n6300), .ZN(n6305) );
  INV_X1 U3466 ( .A(n6300), .ZN(n6306) );
  INV_X1 U3467 ( .A(n6300), .ZN(n6307) );
  INV_X1 U3468 ( .A(n4436), .ZN(n6308) );
  INV_X1 U3469 ( .A(n6308), .ZN(n6309) );
  INV_X1 U3470 ( .A(n6308), .ZN(n6310) );
  INV_X1 U3471 ( .A(n6308), .ZN(n6311) );
  INV_X1 U3472 ( .A(n6308), .ZN(n6312) );
  INV_X1 U3473 ( .A(n6308), .ZN(n6313) );
  INV_X1 U3474 ( .A(n6308), .ZN(n6314) );
  INV_X1 U3475 ( .A(n6308), .ZN(n6315) );
  INV_X1 U3476 ( .A(n4437), .ZN(n6316) );
  INV_X1 U3477 ( .A(n6316), .ZN(n6317) );
  INV_X1 U3478 ( .A(n6316), .ZN(n6318) );
  INV_X1 U3479 ( .A(n6316), .ZN(n6319) );
  INV_X1 U3480 ( .A(n6316), .ZN(n6320) );
  INV_X1 U3481 ( .A(n6316), .ZN(n6321) );
  INV_X1 U3482 ( .A(n6316), .ZN(n6322) );
  INV_X1 U3483 ( .A(n6316), .ZN(n6323) );
  INV_X1 U3484 ( .A(n6324), .ZN(n6325) );
  INV_X1 U3485 ( .A(n6324), .ZN(n6326) );
  INV_X1 U3486 ( .A(n6324), .ZN(n6327) );
  INV_X1 U3487 ( .A(n6324), .ZN(n6328) );
  INV_X1 U3488 ( .A(n6324), .ZN(n6329) );
  INV_X1 U3489 ( .A(n6324), .ZN(n6330) );
  INV_X1 U3490 ( .A(n6324), .ZN(n6331) );
  INV_X1 U3491 ( .A(n4431), .ZN(n6339) );
  INV_X1 U3492 ( .A(n4431), .ZN(n6340) );
  INV_X1 U3493 ( .A(n6339), .ZN(n6341) );
  INV_X1 U3494 ( .A(n6339), .ZN(n6342) );
  INV_X1 U3495 ( .A(n6340), .ZN(n6343) );
  INV_X1 U3496 ( .A(n6339), .ZN(n6344) );
  INV_X1 U3497 ( .A(n6340), .ZN(n6345) );
  INV_X1 U3498 ( .A(n6340), .ZN(n6346) );
  INV_X1 U3499 ( .A(n4432), .ZN(n6347) );
  INV_X1 U3500 ( .A(n6347), .ZN(n6348) );
  INV_X1 U3501 ( .A(n6347), .ZN(n6349) );
  INV_X1 U3502 ( .A(n6347), .ZN(n6350) );
  INV_X1 U3503 ( .A(n6347), .ZN(n6351) );
  INV_X1 U3504 ( .A(n6347), .ZN(n6352) );
  INV_X1 U3505 ( .A(n6347), .ZN(n6353) );
  INV_X1 U3506 ( .A(n6347), .ZN(n6354) );
  INV_X1 U3507 ( .A(n6355), .ZN(n6356) );
  INV_X1 U3508 ( .A(n6355), .ZN(n6357) );
  INV_X1 U3509 ( .A(n6355), .ZN(n6358) );
  INV_X1 U3510 ( .A(n6355), .ZN(n6359) );
  INV_X1 U3511 ( .A(n6355), .ZN(n6360) );
  INV_X1 U3512 ( .A(n6355), .ZN(n6361) );
  INV_X1 U3513 ( .A(n6355), .ZN(n6362) );
  INV_X1 U3514 ( .A(n6363), .ZN(n6364) );
  INV_X1 U3515 ( .A(n6363), .ZN(n6365) );
  INV_X1 U3516 ( .A(n6363), .ZN(n6366) );
  INV_X1 U3517 ( .A(n6363), .ZN(n6367) );
  INV_X1 U3518 ( .A(n6363), .ZN(n6368) );
  INV_X1 U3519 ( .A(n6363), .ZN(n6369) );
  INV_X1 U3520 ( .A(n6363), .ZN(n6370) );
  INV_X1 U3521 ( .A(n4426), .ZN(n6371) );
  INV_X1 U3522 ( .A(n6371), .ZN(n6372) );
  INV_X1 U3523 ( .A(n6371), .ZN(n6373) );
  INV_X1 U3524 ( .A(n6371), .ZN(n6374) );
  INV_X1 U3525 ( .A(n6371), .ZN(n6375) );
  INV_X1 U3526 ( .A(n6371), .ZN(n6376) );
  INV_X1 U3527 ( .A(n6371), .ZN(n6377) );
  INV_X1 U3528 ( .A(n6371), .ZN(n6378) );
  INV_X1 U3529 ( .A(n6395), .ZN(n6396) );
  INV_X1 U3530 ( .A(n6395), .ZN(n6397) );
  INV_X1 U3531 ( .A(n6395), .ZN(n6398) );
  INV_X1 U3532 ( .A(n6395), .ZN(n6399) );
  INV_X1 U3533 ( .A(n6395), .ZN(n6400) );
  INV_X1 U3534 ( .A(n6395), .ZN(n6401) );
  INV_X1 U3535 ( .A(n6395), .ZN(n6402) );
  INV_X1 U3536 ( .A(n6403), .ZN(n6404) );
  INV_X1 U3537 ( .A(n6403), .ZN(n6405) );
  INV_X1 U3538 ( .A(n6403), .ZN(n6406) );
  INV_X1 U3539 ( .A(n6403), .ZN(n6407) );
  INV_X1 U3540 ( .A(n6403), .ZN(n6408) );
  INV_X1 U3541 ( .A(n6403), .ZN(n6409) );
  INV_X1 U3542 ( .A(n6403), .ZN(n6410) );
  INV_X1 U3543 ( .A(n4412), .ZN(n6411) );
  INV_X1 U3544 ( .A(n6411), .ZN(n6412) );
  INV_X1 U3545 ( .A(n6411), .ZN(n6413) );
  INV_X1 U3546 ( .A(n6411), .ZN(n6414) );
  INV_X1 U3547 ( .A(n6411), .ZN(n6415) );
  INV_X1 U3548 ( .A(n6411), .ZN(n6416) );
  INV_X1 U3549 ( .A(n6411), .ZN(n6417) );
  INV_X1 U3550 ( .A(n6411), .ZN(n6418) );
  INV_X1 U3551 ( .A(n4407), .ZN(n6431) );
  INV_X1 U3552 ( .A(n6431), .ZN(n6432) );
  INV_X1 U3553 ( .A(n6431), .ZN(n6433) );
  INV_X1 U3554 ( .A(n6431), .ZN(n6434) );
  INV_X1 U3555 ( .A(n6431), .ZN(n6435) );
  INV_X1 U3556 ( .A(n6431), .ZN(n6436) );
  INV_X1 U3557 ( .A(n6431), .ZN(n6437) );
  INV_X1 U3558 ( .A(n6431), .ZN(n6438) );
  INV_X1 U3559 ( .A(n4408), .ZN(n6439) );
  INV_X1 U3560 ( .A(n6439), .ZN(n6440) );
  INV_X1 U3561 ( .A(n6439), .ZN(n6441) );
  INV_X1 U3562 ( .A(n6439), .ZN(n6442) );
  INV_X1 U3563 ( .A(n6439), .ZN(n6443) );
  INV_X1 U3564 ( .A(n6439), .ZN(n6444) );
  INV_X1 U3565 ( .A(n6439), .ZN(n6445) );
  INV_X1 U3566 ( .A(n6439), .ZN(n6446) );
  INV_X1 U3567 ( .A(n6447), .ZN(n6448) );
  INV_X1 U3568 ( .A(n6447), .ZN(n6449) );
  INV_X1 U3569 ( .A(n6447), .ZN(n6450) );
  INV_X1 U3570 ( .A(n6447), .ZN(n6451) );
  INV_X1 U3571 ( .A(n6447), .ZN(n6452) );
  INV_X1 U3572 ( .A(n6447), .ZN(n6453) );
  INV_X1 U3573 ( .A(n6447), .ZN(n6454) );
  INV_X1 U3574 ( .A(n6455), .ZN(n6456) );
  INV_X1 U3575 ( .A(n6455), .ZN(n6457) );
  INV_X1 U3576 ( .A(n6455), .ZN(n6458) );
  INV_X1 U3577 ( .A(n6455), .ZN(n6459) );
  INV_X1 U3578 ( .A(n6455), .ZN(n6460) );
  INV_X1 U3579 ( .A(n6455), .ZN(n6461) );
  INV_X1 U3580 ( .A(n6455), .ZN(n6462) );
  INV_X1 U3581 ( .A(n6472), .ZN(n6473) );
  INV_X1 U3582 ( .A(n6472), .ZN(n6474) );
  INV_X1 U3583 ( .A(n6472), .ZN(n6475) );
  INV_X1 U3584 ( .A(n6472), .ZN(n6476) );
  INV_X1 U3585 ( .A(n6472), .ZN(n6477) );
  INV_X1 U3586 ( .A(n6472), .ZN(n6478) );
  INV_X1 U3587 ( .A(n6472), .ZN(n6479) );
  INV_X1 U3588 ( .A(n6480), .ZN(n6481) );
  INV_X1 U3589 ( .A(n6480), .ZN(n6482) );
  INV_X1 U3590 ( .A(n6480), .ZN(n6483) );
  INV_X1 U3591 ( .A(n6480), .ZN(n6484) );
  INV_X1 U3592 ( .A(n6480), .ZN(n6485) );
  INV_X1 U3593 ( .A(n6480), .ZN(n6486) );
  INV_X1 U3594 ( .A(n6480), .ZN(n6487) );
  INV_X1 U3595 ( .A(n6491), .ZN(n6493) );
  INV_X1 U3596 ( .A(n6491), .ZN(n6494) );
  INV_X1 U3597 ( .A(n6491), .ZN(n6495) );
  INV_X1 U3598 ( .A(n6492), .ZN(n6496) );
  INV_X1 U3599 ( .A(n6492), .ZN(n6497) );
  INV_X1 U3600 ( .A(n6491), .ZN(n6498) );
  INV_X1 U3601 ( .A(n6491), .ZN(n6499) );
  INV_X1 U3602 ( .A(n6500), .ZN(n6502) );
  INV_X1 U3603 ( .A(n6500), .ZN(n6503) );
  INV_X1 U3604 ( .A(n6500), .ZN(n6504) );
  INV_X1 U3605 ( .A(n6501), .ZN(n6505) );
  INV_X1 U3606 ( .A(n6501), .ZN(n6506) );
  INV_X1 U3607 ( .A(n6500), .ZN(n6507) );
  INV_X1 U3608 ( .A(n6500), .ZN(n6508) );
  INV_X1 U3609 ( .A(n6510), .ZN(n6511) );
  INV_X1 U3610 ( .A(n6509), .ZN(n6512) );
  INV_X1 U3611 ( .A(n6509), .ZN(n6513) );
  INV_X1 U3612 ( .A(n6509), .ZN(n6514) );
  INV_X1 U3613 ( .A(n6510), .ZN(n6515) );
  INV_X1 U3614 ( .A(n6510), .ZN(n6516) );
  INV_X1 U3615 ( .A(n6517), .ZN(n6519) );
  INV_X1 U3616 ( .A(n6517), .ZN(n6520) );
  INV_X1 U3617 ( .A(n6517), .ZN(n6521) );
  INV_X1 U3618 ( .A(n6518), .ZN(n6522) );
  INV_X1 U3619 ( .A(n6518), .ZN(n6523) );
  INV_X1 U3620 ( .A(n6518), .ZN(n6524) );
  INV_X1 U3621 ( .A(n6526), .ZN(n6527) );
  INV_X1 U3622 ( .A(n6525), .ZN(n6528) );
  INV_X1 U3623 ( .A(n6525), .ZN(n6529) );
  INV_X1 U3624 ( .A(n6525), .ZN(n6530) );
  INV_X1 U3625 ( .A(n6526), .ZN(n6531) );
  INV_X1 U3626 ( .A(n6526), .ZN(n6532) );
  INV_X1 U3627 ( .A(n6533), .ZN(n6534) );
  INV_X1 U3628 ( .A(n6533), .ZN(n6535) );
  INV_X1 U3629 ( .A(n6533), .ZN(n6536) );
  INV_X1 U3630 ( .A(n6533), .ZN(n6537) );
  INV_X1 U3631 ( .A(n6533), .ZN(n6538) );
  INV_X1 U3632 ( .A(n6533), .ZN(n6539) );
  INV_X1 U3633 ( .A(n6533), .ZN(n6540) );
  INV_X1 U3634 ( .A(n6533), .ZN(n6541) );
  INV_X1 U3635 ( .A(n6543), .ZN(n6544) );
  INV_X1 U3636 ( .A(n6542), .ZN(n6545) );
  INV_X1 U3637 ( .A(n6542), .ZN(n6546) );
  INV_X1 U3638 ( .A(n6542), .ZN(n6547) );
  INV_X1 U3639 ( .A(n6543), .ZN(n6548) );
  INV_X1 U3640 ( .A(n6543), .ZN(n6549) );
  INV_X1 U3641 ( .A(n6550), .ZN(n6552) );
  INV_X1 U3642 ( .A(n6550), .ZN(n6553) );
  INV_X1 U3643 ( .A(n6550), .ZN(n6554) );
  INV_X1 U3644 ( .A(n6551), .ZN(n6555) );
  INV_X1 U3645 ( .A(n6551), .ZN(n6556) );
  INV_X1 U3646 ( .A(n6551), .ZN(n6557) );
  INV_X1 U3647 ( .A(n6558), .ZN(n6560) );
  INV_X1 U3648 ( .A(n6558), .ZN(n6561) );
  INV_X1 U3649 ( .A(n6558), .ZN(n6562) );
  INV_X1 U3650 ( .A(n6559), .ZN(n6563) );
  INV_X1 U3651 ( .A(n6559), .ZN(n6564) );
  INV_X1 U3652 ( .A(n6558), .ZN(n6565) );
  INV_X1 U3653 ( .A(n6558), .ZN(n6566) );
  INV_X1 U3654 ( .A(n6567), .ZN(n6569) );
  INV_X1 U3655 ( .A(n6567), .ZN(n6570) );
  INV_X1 U3656 ( .A(n6567), .ZN(n6571) );
  INV_X1 U3657 ( .A(n6568), .ZN(n6572) );
  INV_X1 U3658 ( .A(n6568), .ZN(n6573) );
  INV_X1 U3659 ( .A(n6567), .ZN(n6574) );
  INV_X1 U3660 ( .A(n6567), .ZN(n6575) );
  INV_X1 U3661 ( .A(n6576), .ZN(n6578) );
  INV_X1 U3662 ( .A(n6576), .ZN(n6579) );
  INV_X1 U3663 ( .A(n6576), .ZN(n6580) );
  INV_X1 U3664 ( .A(n6577), .ZN(n6581) );
  INV_X1 U3665 ( .A(n6577), .ZN(n6582) );
  INV_X1 U3666 ( .A(n6576), .ZN(n6583) );
  INV_X1 U3667 ( .A(n6576), .ZN(n6584) );
  INV_X1 U3668 ( .A(n6585), .ZN(n6587) );
  INV_X1 U3669 ( .A(n6585), .ZN(n6588) );
  INV_X1 U3670 ( .A(n6585), .ZN(n6589) );
  INV_X1 U3671 ( .A(n6586), .ZN(n6590) );
  INV_X1 U3672 ( .A(n6586), .ZN(n6591) );
  INV_X1 U3673 ( .A(n6585), .ZN(n6592) );
  INV_X1 U3674 ( .A(n6585), .ZN(n6593) );
  INV_X1 U3675 ( .A(n6595), .ZN(n6596) );
  INV_X1 U3676 ( .A(n6594), .ZN(n6597) );
  INV_X1 U3677 ( .A(n6594), .ZN(n6598) );
  INV_X1 U3678 ( .A(n6594), .ZN(n6599) );
  INV_X1 U3679 ( .A(n6595), .ZN(n6600) );
  INV_X1 U3680 ( .A(n6595), .ZN(n6601) );
  INV_X1 U3681 ( .A(n6602), .ZN(n6603) );
  INV_X1 U3682 ( .A(n6602), .ZN(n6604) );
  INV_X1 U3683 ( .A(n6602), .ZN(n6605) );
  INV_X1 U3684 ( .A(n6602), .ZN(n6606) );
  INV_X1 U3685 ( .A(n6602), .ZN(n6607) );
  INV_X1 U3686 ( .A(n6602), .ZN(n6608) );
  INV_X1 U3687 ( .A(n6602), .ZN(n6609) );
  INV_X1 U3688 ( .A(n6602), .ZN(n6610) );
  INV_X1 U3689 ( .A(n6612), .ZN(n6613) );
  INV_X1 U3690 ( .A(n6611), .ZN(n6614) );
  INV_X1 U3691 ( .A(n6611), .ZN(n6615) );
  INV_X1 U3692 ( .A(n6611), .ZN(n6616) );
  INV_X1 U3693 ( .A(n6612), .ZN(n6617) );
  INV_X1 U3694 ( .A(n6612), .ZN(n6618) );
  INV_X1 U3695 ( .A(n6619), .ZN(n6621) );
  INV_X1 U3696 ( .A(n6619), .ZN(n6622) );
  INV_X1 U3697 ( .A(n6619), .ZN(n6623) );
  INV_X1 U3698 ( .A(n6620), .ZN(n6624) );
  INV_X1 U3699 ( .A(n6620), .ZN(n6625) );
  INV_X1 U3700 ( .A(n6620), .ZN(n6626) );
  INV_X1 U3701 ( .A(n6627), .ZN(n6629) );
  INV_X1 U3702 ( .A(n6627), .ZN(n6630) );
  INV_X1 U3703 ( .A(n6627), .ZN(n6631) );
  INV_X1 U3704 ( .A(n6628), .ZN(n6632) );
  INV_X1 U3705 ( .A(n6628), .ZN(n6633) );
  INV_X1 U3706 ( .A(n6627), .ZN(n6634) );
  INV_X1 U3707 ( .A(n6627), .ZN(n6635) );
  INV_X1 U3708 ( .A(n6636), .ZN(n6638) );
  INV_X1 U3709 ( .A(n6636), .ZN(n6639) );
  INV_X1 U3710 ( .A(n6636), .ZN(n6640) );
  INV_X1 U3711 ( .A(n6637), .ZN(n6641) );
  INV_X1 U3712 ( .A(n6637), .ZN(n6642) );
  INV_X1 U3713 ( .A(n6636), .ZN(n6643) );
  INV_X1 U3714 ( .A(n6636), .ZN(n6644) );
  INV_X1 U3715 ( .A(n6645), .ZN(n6647) );
  INV_X1 U3716 ( .A(n6645), .ZN(n6648) );
  INV_X1 U3717 ( .A(n6645), .ZN(n6649) );
  INV_X1 U3718 ( .A(n6646), .ZN(n6650) );
  INV_X1 U3719 ( .A(n6646), .ZN(n6651) );
  INV_X1 U3720 ( .A(n6645), .ZN(n6652) );
  INV_X1 U3721 ( .A(n6645), .ZN(n6653) );
  INV_X1 U3722 ( .A(n6654), .ZN(n6656) );
  INV_X1 U3723 ( .A(n6654), .ZN(n6657) );
  INV_X1 U3724 ( .A(n6654), .ZN(n6658) );
  INV_X1 U3725 ( .A(n6655), .ZN(n6659) );
  INV_X1 U3726 ( .A(n6655), .ZN(n6660) );
  INV_X1 U3727 ( .A(n6654), .ZN(n6661) );
  INV_X1 U3728 ( .A(n6654), .ZN(n6662) );
  INV_X1 U3729 ( .A(n6663), .ZN(n6665) );
  INV_X1 U3730 ( .A(n6663), .ZN(n6666) );
  INV_X1 U3731 ( .A(n6663), .ZN(n6667) );
  INV_X1 U3732 ( .A(n6663), .ZN(n6668) );
  INV_X1 U3733 ( .A(n6663), .ZN(n6669) );
  INV_X1 U3734 ( .A(n6663), .ZN(n6670) );
  INV_X1 U3735 ( .A(n6664), .ZN(n6671) );
  INV_X1 U3736 ( .A(n6673), .ZN(n6674) );
  INV_X1 U3737 ( .A(n6672), .ZN(n6675) );
  INV_X1 U3738 ( .A(n6672), .ZN(n6676) );
  INV_X1 U3739 ( .A(n6673), .ZN(n6677) );
  INV_X1 U3740 ( .A(n6673), .ZN(n6678) );
  INV_X1 U3741 ( .A(n6673), .ZN(n6679) );
  INV_X1 U3742 ( .A(n6673), .ZN(n6680) );
  INV_X1 U3743 ( .A(n6681), .ZN(n6683) );
  INV_X1 U3744 ( .A(n6681), .ZN(n6684) );
  INV_X1 U3745 ( .A(n6681), .ZN(n6685) );
  INV_X1 U3746 ( .A(n6681), .ZN(n6686) );
  INV_X1 U3747 ( .A(n6681), .ZN(n6687) );
  INV_X1 U3748 ( .A(n6681), .ZN(n6688) );
  INV_X1 U3749 ( .A(n6682), .ZN(n6689) );
  INV_X1 U3750 ( .A(n6691), .ZN(n6692) );
  INV_X1 U3751 ( .A(n6690), .ZN(n6693) );
  INV_X1 U3752 ( .A(n6690), .ZN(n6694) );
  INV_X1 U3753 ( .A(n6691), .ZN(n6695) );
  INV_X1 U3754 ( .A(n6691), .ZN(n6696) );
  INV_X1 U3755 ( .A(n6691), .ZN(n6697) );
  INV_X1 U3756 ( .A(n6691), .ZN(n6698) );
  INV_X1 U3757 ( .A(n6713), .ZN(n6715) );
  INV_X1 U3758 ( .A(n6713), .ZN(n6716) );
  INV_X1 U3759 ( .A(n6713), .ZN(n6717) );
  INV_X1 U3760 ( .A(n6714), .ZN(n6718) );
  INV_X1 U3761 ( .A(n6714), .ZN(n6719) );
  INV_X1 U3762 ( .A(n6713), .ZN(n6720) );
  INV_X1 U3763 ( .A(n6713), .ZN(n6721) );
  INV_X1 U3764 ( .A(n6722), .ZN(n6724) );
  INV_X1 U3765 ( .A(n6722), .ZN(n6725) );
  INV_X1 U3766 ( .A(n6722), .ZN(n6726) );
  INV_X1 U3767 ( .A(n6723), .ZN(n6727) );
  INV_X1 U3768 ( .A(n6723), .ZN(n6728) );
  INV_X1 U3769 ( .A(n6722), .ZN(n6729) );
  INV_X1 U3770 ( .A(n6722), .ZN(n6730) );
  CLKBUF_X1 U3771 ( .A(n6872), .Z(n6766) );
  CLKBUF_X1 U3772 ( .A(n6871), .Z(n6767) );
  CLKBUF_X1 U3773 ( .A(n6871), .Z(n6768) );
  CLKBUF_X1 U3774 ( .A(n6871), .Z(n6769) );
  CLKBUF_X1 U3775 ( .A(n6871), .Z(n6770) );
  CLKBUF_X1 U3776 ( .A(n6871), .Z(n6771) );
  CLKBUF_X1 U3777 ( .A(n6871), .Z(n6772) );
  CLKBUF_X1 U3778 ( .A(n6870), .Z(n6773) );
  CLKBUF_X1 U3779 ( .A(n6870), .Z(n6774) );
  CLKBUF_X1 U3780 ( .A(n6870), .Z(n6775) );
  CLKBUF_X1 U3781 ( .A(n6870), .Z(n6776) );
  CLKBUF_X1 U3782 ( .A(n6870), .Z(n6777) );
  CLKBUF_X1 U3783 ( .A(n6870), .Z(n6778) );
  CLKBUF_X1 U3784 ( .A(n6869), .Z(n6779) );
  CLKBUF_X1 U3785 ( .A(n6869), .Z(n6780) );
  CLKBUF_X1 U3786 ( .A(n6869), .Z(n6781) );
  CLKBUF_X1 U3787 ( .A(n6869), .Z(n6782) );
  CLKBUF_X1 U3788 ( .A(n6869), .Z(n6783) );
  CLKBUF_X1 U3789 ( .A(n6869), .Z(n6784) );
  CLKBUF_X1 U3790 ( .A(n6868), .Z(n6785) );
  CLKBUF_X1 U3791 ( .A(n6868), .Z(n6786) );
  CLKBUF_X1 U3792 ( .A(n6868), .Z(n6787) );
  CLKBUF_X1 U3793 ( .A(n6868), .Z(n6788) );
  CLKBUF_X1 U3794 ( .A(n6868), .Z(n6789) );
  CLKBUF_X1 U3795 ( .A(n6868), .Z(n6790) );
  CLKBUF_X1 U3796 ( .A(n6867), .Z(n6791) );
  CLKBUF_X1 U3797 ( .A(n6867), .Z(n6792) );
  CLKBUF_X1 U3798 ( .A(n6867), .Z(n6793) );
  CLKBUF_X1 U3799 ( .A(n6867), .Z(n6794) );
  CLKBUF_X1 U3800 ( .A(n6867), .Z(n6795) );
  CLKBUF_X1 U3801 ( .A(n6867), .Z(n6796) );
  CLKBUF_X1 U3802 ( .A(n6866), .Z(n6797) );
  CLKBUF_X1 U3803 ( .A(n6866), .Z(n6798) );
  CLKBUF_X1 U3804 ( .A(n6866), .Z(n6799) );
  CLKBUF_X1 U3805 ( .A(n6866), .Z(n6800) );
  CLKBUF_X1 U3806 ( .A(n6866), .Z(n6801) );
  CLKBUF_X1 U3807 ( .A(n6866), .Z(n6802) );
  CLKBUF_X1 U3808 ( .A(n6865), .Z(n6803) );
  CLKBUF_X1 U3809 ( .A(n6865), .Z(n6804) );
  CLKBUF_X1 U3810 ( .A(n6865), .Z(n6805) );
  CLKBUF_X1 U3811 ( .A(n6865), .Z(n6806) );
  CLKBUF_X1 U3812 ( .A(n6865), .Z(n6807) );
  CLKBUF_X1 U3813 ( .A(n6865), .Z(n6808) );
  CLKBUF_X1 U3814 ( .A(n6864), .Z(n6809) );
  CLKBUF_X1 U3815 ( .A(n6864), .Z(n6810) );
  CLKBUF_X1 U3816 ( .A(n6864), .Z(n6811) );
  CLKBUF_X1 U3817 ( .A(n6864), .Z(n6812) );
  CLKBUF_X1 U3818 ( .A(n6864), .Z(n6813) );
  CLKBUF_X1 U3819 ( .A(n6864), .Z(n6814) );
  CLKBUF_X1 U3820 ( .A(n6863), .Z(n6815) );
  CLKBUF_X1 U3821 ( .A(n6863), .Z(n6816) );
  CLKBUF_X1 U3822 ( .A(n6863), .Z(n6817) );
  CLKBUF_X1 U3823 ( .A(n6863), .Z(n6818) );
  CLKBUF_X1 U3824 ( .A(n6863), .Z(n6819) );
  CLKBUF_X1 U3825 ( .A(n6863), .Z(n6820) );
  CLKBUF_X1 U3826 ( .A(n6862), .Z(n6821) );
  CLKBUF_X1 U3827 ( .A(n6862), .Z(n6822) );
  CLKBUF_X1 U3828 ( .A(n6862), .Z(n6823) );
  CLKBUF_X1 U3829 ( .A(n6862), .Z(n6824) );
  CLKBUF_X1 U3830 ( .A(n6862), .Z(n6825) );
  CLKBUF_X1 U3831 ( .A(n6862), .Z(n6826) );
  CLKBUF_X1 U3832 ( .A(n6861), .Z(n6827) );
  CLKBUF_X1 U3833 ( .A(n6861), .Z(n6828) );
  CLKBUF_X1 U3834 ( .A(n6861), .Z(n6829) );
  CLKBUF_X1 U3835 ( .A(n6861), .Z(n6830) );
  CLKBUF_X1 U3836 ( .A(n6861), .Z(n6831) );
  CLKBUF_X1 U3837 ( .A(n6861), .Z(n6832) );
  CLKBUF_X1 U3838 ( .A(n6860), .Z(n6833) );
  CLKBUF_X1 U3839 ( .A(n6860), .Z(n6834) );
  CLKBUF_X1 U3840 ( .A(n6860), .Z(n6835) );
  CLKBUF_X1 U3841 ( .A(n6860), .Z(n6836) );
  CLKBUF_X1 U3842 ( .A(n6860), .Z(n6837) );
  CLKBUF_X1 U3843 ( .A(n6860), .Z(n6838) );
  CLKBUF_X1 U3844 ( .A(n6859), .Z(n6839) );
  CLKBUF_X1 U3845 ( .A(n6859), .Z(n6840) );
  CLKBUF_X1 U3846 ( .A(n6859), .Z(n6841) );
  CLKBUF_X1 U3847 ( .A(n6859), .Z(n6842) );
  CLKBUF_X1 U3848 ( .A(n6859), .Z(n6843) );
  CLKBUF_X1 U3849 ( .A(n6859), .Z(n6844) );
  CLKBUF_X1 U3850 ( .A(n6858), .Z(n6845) );
  CLKBUF_X1 U3851 ( .A(n6858), .Z(n6846) );
  CLKBUF_X1 U3852 ( .A(n6858), .Z(n6847) );
  CLKBUF_X1 U3853 ( .A(n6858), .Z(n6848) );
  CLKBUF_X1 U3854 ( .A(n6858), .Z(n6849) );
  CLKBUF_X1 U3855 ( .A(n6858), .Z(n6850) );
  CLKBUF_X1 U3856 ( .A(n6857), .Z(n6851) );
  CLKBUF_X1 U3857 ( .A(n6857), .Z(n6852) );
  CLKBUF_X1 U3858 ( .A(n6857), .Z(n6853) );
  CLKBUF_X1 U3859 ( .A(n6857), .Z(n6854) );
  CLKBUF_X1 U3860 ( .A(n6857), .Z(n6855) );
  CLKBUF_X1 U3861 ( .A(n6857), .Z(n6856) );
endmodule


module rca_n_n32_0 ( a, b, c_in, sum, c_out );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input c_in;
  output c_out;

  wire   [31:1] temp;

  fa_2_0 fa_2_i_0 ( .a(a[0]), .b(b[0]), .c_in(c_in), .sum(sum[0]), .c_out(
        temp[1]) );
  fa_2_159 fa_2_i_1 ( .a(a[1]), .b(b[1]), .c_in(temp[1]), .sum(sum[1]), 
        .c_out(temp[2]) );
  fa_2_158 fa_2_i_2 ( .a(a[2]), .b(b[2]), .c_in(temp[2]), .sum(sum[2]), 
        .c_out(temp[3]) );
  fa_2_157 fa_2_i_3 ( .a(a[3]), .b(b[3]), .c_in(temp[3]), .sum(sum[3]), 
        .c_out(temp[4]) );
  fa_2_156 fa_2_i_4 ( .a(a[4]), .b(b[4]), .c_in(temp[4]), .sum(sum[4]), 
        .c_out(temp[5]) );
  fa_2_155 fa_2_i_5 ( .a(a[5]), .b(b[5]), .c_in(temp[5]), .sum(sum[5]), 
        .c_out(temp[6]) );
  fa_2_154 fa_2_i_6 ( .a(a[6]), .b(b[6]), .c_in(temp[6]), .sum(sum[6]), 
        .c_out(temp[7]) );
  fa_2_153 fa_2_i_7 ( .a(a[7]), .b(b[7]), .c_in(temp[7]), .sum(sum[7]), 
        .c_out(temp[8]) );
  fa_2_152 fa_2_i_8 ( .a(a[8]), .b(b[8]), .c_in(temp[8]), .sum(sum[8]), 
        .c_out(temp[9]) );
  fa_2_151 fa_2_i_9 ( .a(a[9]), .b(b[9]), .c_in(temp[9]), .sum(sum[9]), 
        .c_out(temp[10]) );
  fa_2_150 fa_2_i_10 ( .a(a[10]), .b(b[10]), .c_in(temp[10]), .sum(sum[10]), 
        .c_out(temp[11]) );
  fa_2_149 fa_2_i_11 ( .a(a[11]), .b(b[11]), .c_in(temp[11]), .sum(sum[11]), 
        .c_out(temp[12]) );
  fa_2_148 fa_2_i_12 ( .a(a[12]), .b(b[12]), .c_in(temp[12]), .sum(sum[12]), 
        .c_out(temp[13]) );
  fa_2_147 fa_2_i_13 ( .a(a[13]), .b(b[13]), .c_in(temp[13]), .sum(sum[13]), 
        .c_out(temp[14]) );
  fa_2_146 fa_2_i_14 ( .a(a[14]), .b(b[14]), .c_in(temp[14]), .sum(sum[14]), 
        .c_out(temp[15]) );
  fa_2_145 fa_2_i_15 ( .a(a[15]), .b(b[15]), .c_in(temp[15]), .sum(sum[15]), 
        .c_out(temp[16]) );
  fa_2_144 fa_2_i_16 ( .a(a[16]), .b(b[16]), .c_in(temp[16]), .sum(sum[16]), 
        .c_out(temp[17]) );
  fa_2_143 fa_2_i_17 ( .a(a[17]), .b(b[17]), .c_in(temp[17]), .sum(sum[17]), 
        .c_out(temp[18]) );
  fa_2_142 fa_2_i_18 ( .a(a[18]), .b(b[18]), .c_in(temp[18]), .sum(sum[18]), 
        .c_out(temp[19]) );
  fa_2_141 fa_2_i_19 ( .a(a[19]), .b(b[19]), .c_in(temp[19]), .sum(sum[19]), 
        .c_out(temp[20]) );
  fa_2_140 fa_2_i_20 ( .a(a[20]), .b(b[20]), .c_in(temp[20]), .sum(sum[20]), 
        .c_out(temp[21]) );
  fa_2_139 fa_2_i_21 ( .a(a[21]), .b(b[21]), .c_in(temp[21]), .sum(sum[21]), 
        .c_out(temp[22]) );
  fa_2_138 fa_2_i_22 ( .a(a[22]), .b(b[22]), .c_in(temp[22]), .sum(sum[22]), 
        .c_out(temp[23]) );
  fa_2_137 fa_2_i_23 ( .a(a[23]), .b(b[23]), .c_in(temp[23]), .sum(sum[23]), 
        .c_out(temp[24]) );
  fa_2_136 fa_2_i_24 ( .a(a[24]), .b(b[24]), .c_in(temp[24]), .sum(sum[24]), 
        .c_out(temp[25]) );
  fa_2_135 fa_2_i_25 ( .a(a[25]), .b(b[25]), .c_in(temp[25]), .sum(sum[25]), 
        .c_out(temp[26]) );
  fa_2_134 fa_2_i_26 ( .a(a[26]), .b(b[26]), .c_in(temp[26]), .sum(sum[26]), 
        .c_out(temp[27]) );
  fa_2_133 fa_2_i_27 ( .a(a[27]), .b(b[27]), .c_in(temp[27]), .sum(sum[27]), 
        .c_out(temp[28]) );
  fa_2_132 fa_2_i_28 ( .a(a[28]), .b(b[28]), .c_in(temp[28]), .sum(sum[28]), 
        .c_out(temp[29]) );
  fa_2_131 fa_2_i_29 ( .a(a[29]), .b(b[29]), .c_in(temp[29]), .sum(sum[29]), 
        .c_out(temp[30]) );
  fa_2_130 fa_2_i_30 ( .a(a[30]), .b(b[30]), .c_in(temp[30]), .sum(sum[30]), 
        .c_out(temp[31]) );
  fa_2_129 fa_2_i_31 ( .a(a[31]), .b(b[31]), .c_in(temp[31]), .sum(sum[31]), 
        .c_out(c_out) );
endmodule


module reg_n_n32_0 ( clock, reset, enable, x, y );
  input [31:0] x;
  output [31:0] y;
  input clock, reset, enable;
  wire   n1, n2, n3;

  ffd_async_271 ff_0 ( .clk(clock), .reset(n1), .en(enable), .d(x[0]), .q(y[0]) );
  ffd_async_270 ff_1 ( .clk(clock), .reset(n1), .en(enable), .d(x[1]), .q(y[1]) );
  ffd_async_269 ff_2 ( .clk(clock), .reset(n1), .en(enable), .d(x[2]), .q(y[2]) );
  ffd_async_268 ff_3 ( .clk(clock), .reset(n1), .en(enable), .d(x[3]), .q(y[3]) );
  ffd_async_267 ff_4 ( .clk(clock), .reset(n1), .en(enable), .d(x[4]), .q(y[4]) );
  ffd_async_266 ff_5 ( .clk(clock), .reset(n1), .en(enable), .d(x[5]), .q(y[5]) );
  ffd_async_265 ff_6 ( .clk(clock), .reset(n1), .en(enable), .d(x[6]), .q(y[6]) );
  ffd_async_264 ff_7 ( .clk(clock), .reset(n1), .en(enable), .d(x[7]), .q(y[7]) );
  ffd_async_263 ff_8 ( .clk(clock), .reset(n1), .en(enable), .d(x[8]), .q(y[8]) );
  ffd_async_262 ff_9 ( .clk(clock), .reset(n1), .en(enable), .d(x[9]), .q(y[9]) );
  ffd_async_261 ff_10 ( .clk(clock), .reset(n1), .en(enable), .d(x[10]), .q(
        y[10]) );
  ffd_async_260 ff_11 ( .clk(clock), .reset(n1), .en(enable), .d(x[11]), .q(
        y[11]) );
  ffd_async_259 ff_12 ( .clk(clock), .reset(n2), .en(enable), .d(x[12]), .q(
        y[12]) );
  ffd_async_258 ff_13 ( .clk(clock), .reset(n2), .en(enable), .d(x[13]), .q(
        y[13]) );
  ffd_async_257 ff_14 ( .clk(clock), .reset(n2), .en(enable), .d(x[14]), .q(
        y[14]) );
  ffd_async_256 ff_15 ( .clk(clock), .reset(n2), .en(enable), .d(x[15]), .q(
        y[15]) );
  ffd_async_255 ff_16 ( .clk(clock), .reset(n2), .en(enable), .d(x[16]), .q(
        y[16]) );
  ffd_async_254 ff_17 ( .clk(clock), .reset(n2), .en(enable), .d(x[17]), .q(
        y[17]) );
  ffd_async_253 ff_18 ( .clk(clock), .reset(n2), .en(enable), .d(x[18]), .q(
        y[18]) );
  ffd_async_252 ff_19 ( .clk(clock), .reset(n2), .en(enable), .d(x[19]), .q(
        y[19]) );
  ffd_async_251 ff_20 ( .clk(clock), .reset(n2), .en(enable), .d(x[20]), .q(
        y[20]) );
  ffd_async_250 ff_21 ( .clk(clock), .reset(n2), .en(enable), .d(x[21]), .q(
        y[21]) );
  ffd_async_249 ff_22 ( .clk(clock), .reset(n2), .en(enable), .d(x[22]), .q(
        y[22]) );
  ffd_async_248 ff_23 ( .clk(clock), .reset(n2), .en(enable), .d(x[23]), .q(
        y[23]) );
  ffd_async_247 ff_24 ( .clk(clock), .reset(n3), .en(enable), .d(x[24]), .q(
        y[24]) );
  ffd_async_246 ff_25 ( .clk(clock), .reset(n3), .en(enable), .d(x[25]), .q(
        y[25]) );
  ffd_async_245 ff_26 ( .clk(clock), .reset(n3), .en(enable), .d(x[26]), .q(
        y[26]) );
  ffd_async_244 ff_27 ( .clk(clock), .reset(n3), .en(enable), .d(x[27]), .q(
        y[27]) );
  ffd_async_243 ff_28 ( .clk(clock), .reset(n3), .en(enable), .d(x[28]), .q(
        y[28]) );
  ffd_async_242 ff_29 ( .clk(clock), .reset(n3), .en(enable), .d(x[29]), .q(
        y[29]) );
  ffd_async_241 ff_30 ( .clk(clock), .reset(n3), .en(enable), .d(x[30]), .q(
        y[30]) );
  ffd_async_240 ff_31 ( .clk(clock), .reset(n3), .en(enable), .d(x[31]), .q(
        y[31]) );
  BUF_X1 U1 ( .A(reset), .Z(n1) );
  BUF_X1 U2 ( .A(reset), .Z(n2) );
  BUF_X1 U3 ( .A(reset), .Z(n3) );
endmodule


module datapath ( clk, rst, en0, ir, pc_in, en1, rf1, rf2, en2, s1, s2, alu1, 
        alu2, alu3, alu4, eq_cond, jump_en, en3, rw, den, dram_data_in, 
        dram_rw_en, dram_enable, dram_data_out, dram_addr, pc_out, s3, wf1 );
  input [31:0] ir;
  input [31:0] pc_in;
  input [31:0] dram_data_in;
  output [31:0] dram_data_out;
  output [31:0] dram_addr;
  output [31:0] pc_out;
  input clk, rst, en0, en1, rf1, rf2, en2, s1, s2, alu1, alu2, alu3, alu4,
         eq_cond, jump_en, en3, rw, den, s3, wf1;
  output dram_rw_en, dram_enable;
  wire   wf1_st4, z, eq_cond_st2, cond_xor, jump_en_st2, cond, s1_st2, s2_st2,
         en2_st2, en3_st3, s3_st4, en2_st1, s1_st1, s2_st1, alu1_st1, alu2_st1,
         alu3_st1, alu4_st1, eq_cond_st1, jump_en_st1, en3_st1, rw_st1,
         den_st1, s3_st1, wf1_st1, en3_st2, rw_st2, den_st2, s3_st2, wf1_st2,
         s3_st3, wf1_st3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33;
  wire   [31:0] ir_st1;
  wire   [31:0] npc;
  wire   [4:0] rd2;
  wire   [4:0] rd;
  wire   [15:0] inp2;
  wire   [4:0] out_rd3;
  wire   [31:0] wb;
  wire   [31:0] rf_out1;
  wire   [31:0] rf_out2;
  wire   [31:0] out_a;
  wire   [31:0] out_b;
  wire   [31:0] inp2_32;
  wire   [31:0] imm_st2;
  wire   [4:0] out_rd1;
  wire   [3:0] alu_bit;
  wire   [31:0] out_mux1;
  wire   [31:0] out_mux2;
  wire   [31:0] out_alu;
  wire   [4:0] out_rd2;
  wire   [31:0] alu_st4;
  wire   [31:0] out_dram;

  reg_n_n32_0 ir_ff ( .clock(clk), .reset(n32), .enable(en0), .x(ir), .y(
        ir_st1) );
  rca_n_n32_0 pc_add ( .a(pc_in), .b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1}), .c_in(1'b0), .sum(npc) );
  register_file_n32 rf ( .clk(clk), .reset(n32), .enable(en1), .rd1(rf1), 
        .rd2(rf2), .wr(wf1_st4), .add_wr(out_rd3), .add_rd1(ir_st1[25:21]), 
        .add_rd2(rd2), .datain(wb), .out1(rf_out1), .out2(rf_out2) );
  reg_n_n32_7 a ( .clock(clk), .reset(n32), .enable(en1), .x(rf_out1), .y(
        out_a) );
  reg_n_n32_6 b ( .clock(clk), .reset(n32), .enable(en1), .x(rf_out2), .y(
        out_b) );
  sign_extension_s16_f32 ext ( .x(inp2), .y(inp2_32) );
  reg_n_n32_5 in2 ( .clock(clk), .reset(n32), .enable(1'b0), .x(inp2_32), .y(
        imm_st2) );
  reg_n_n5_0 rd_1 ( .clock(clk), .reset(n32), .enable(1'b0), .x(rd), .y(
        out_rd1) );
  zero_comp_n32 cmp ( .x(out_a), .y(z) );
  xor_2_0 eq_xor ( .a(z), .b(eq_cond_st2), .y(cond_xor) );
  and_2_0 and_j ( .a(cond_xor), .b(jump_en_st2), .y(cond) );
  mux21_generic_n32_0 mux1_alu ( .a(npc), .b(out_a), .sel(s1_st2), .y(out_mux1) );
  mux21_generic_n32_3 mux2_alu ( .a(out_b), .b(imm_st2), .sel(s2_st2), .y(
        out_mux2) );
  alu_nbit32 arith_log_un ( .a(out_mux1), .b(out_mux2), .unit_sel(alu_bit), 
        .y(out_alu) );
  reg_n_n32_4 alu_out ( .clock(clk), .reset(n32), .enable(en2_st2), .x(out_alu), .y(dram_addr) );
  reg_n_n32_3 me ( .clock(clk), .reset(n32), .enable(en2_st2), .x(out_b), .y(
        dram_data_out) );
  reg_n_n5_2 rd_2 ( .clock(clk), .reset(n32), .enable(en2_st2), .x(out_rd1), 
        .y(out_rd2) );
  mux21_generic_n32_2 mux_j ( .a(npc), .b(dram_addr), .sel(cond), .y(pc_out)
         );
  reg_n_n32_2 out_value ( .clock(clk), .reset(n32), .enable(en3_st3), .x(
        dram_addr), .y(alu_st4) );
  reg_n_n32_1 lmd ( .clock(clk), .reset(n32), .enable(en3_st3), .x(
        dram_data_in), .y(out_dram) );
  reg_n_n5_1 rd_3 ( .clock(clk), .reset(n32), .enable(en3_st3), .x(out_rd2), 
        .y(out_rd3) );
  mux21_generic_n32_1 mux_out_sel ( .a(out_dram), .b(alu_st4), .sel(s3_st4), 
        .y(wb) );
  ffd_async_0 en2_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(en2), .q(en2_st1) );
  ffd_async_305 s1_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(s1), .q(s1_st1)
         );
  ffd_async_304 s2_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(s2), .q(s2_st1)
         );
  ffd_async_303 alu1_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(alu1), .q(
        alu1_st1) );
  ffd_async_302 alu2_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(alu2), .q(
        alu2_st1) );
  ffd_async_301 alu3_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(alu3), .q(
        alu3_st1) );
  ffd_async_300 alu4_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(alu4), .q(
        alu4_st1) );
  ffd_async_299 eq_cond_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(eq_cond), 
        .q(eq_cond_st1) );
  ffd_async_298 jump_en_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(jump_en), 
        .q(jump_en_st1) );
  ffd_async_297 en3_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(en3), .q(
        en3_st1) );
  ffd_async_296 rw_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(rw), .q(rw_st1)
         );
  ffd_async_295 den_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(den), .q(
        den_st1) );
  ffd_async_294 s3_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(s3), .q(s3_st1)
         );
  ffd_async_293 wf1_cw1 ( .clk(clk), .reset(n33), .en(1'b1), .d(wf1), .q(
        wf1_st1) );
  ffd_async_292 en2_cw2 ( .clk(clk), .reset(n33), .en(1'b1), .d(en2_st1), .q(
        en2_st2) );
  ffd_async_291 s1_cw2 ( .clk(clk), .reset(n33), .en(1'b1), .d(s1_st1), .q(
        s1_st2) );
  ffd_async_290 s2_cw2 ( .clk(clk), .reset(n32), .en(1'b1), .d(s2_st1), .q(
        s2_st2) );
  ffd_async_289 alu1_cw2 ( .clk(clk), .reset(n32), .en(1'b1), .d(alu1_st1), 
        .q(alu_bit[3]) );
  ffd_async_288 alu2_cw2 ( .clk(clk), .reset(n32), .en(1'b1), .d(alu2_st1), 
        .q(alu_bit[2]) );
  ffd_async_287 alu3_cw2 ( .clk(clk), .reset(n32), .en(1'b1), .d(alu3_st1), 
        .q(alu_bit[1]) );
  ffd_async_286 alu4_cw2 ( .clk(clk), .reset(n32), .en(1'b1), .d(alu4_st1), 
        .q(alu_bit[0]) );
  ffd_async_285 eq_cond_cw2 ( .clk(clk), .reset(n33), .en(1'b1), .d(
        eq_cond_st1), .q(eq_cond_st2) );
  ffd_async_284 jump_en_cw2 ( .clk(clk), .reset(n33), .en(1'b1), .d(
        jump_en_st1), .q(jump_en_st2) );
  ffd_async_283 en3_cw2 ( .clk(clk), .reset(n33), .en(1'b1), .d(en3_st1), .q(
        en3_st2) );
  ffd_async_282 rw_cw2 ( .clk(clk), .reset(n33), .en(1'b1), .d(rw_st1), .q(
        rw_st2) );
  ffd_async_281 den_cw2 ( .clk(clk), .reset(n33), .en(1'b1), .d(den_st1), .q(
        den_st2) );
  ffd_async_280 s3_cw2 ( .clk(clk), .reset(n33), .en(1'b1), .d(s3_st1), .q(
        s3_st2) );
  ffd_async_279 wf1_cw2 ( .clk(clk), .reset(n33), .en(1'b1), .d(wf1_st1), .q(
        wf1_st2) );
  ffd_async_278 en3_cw3 ( .clk(clk), .reset(n33), .en(1'b1), .d(en3_st2), .q(
        en3_st3) );
  ffd_async_277 rw_cw3 ( .clk(clk), .reset(n33), .en(1'b1), .d(rw_st2), .q(
        dram_rw_en) );
  ffd_async_276 den_cw3 ( .clk(clk), .reset(n33), .en(1'b1), .d(den_st2), .q(
        dram_enable) );
  ffd_async_275 s3_cw3 ( .clk(clk), .reset(n33), .en(1'b1), .d(s3_st2), .q(
        s3_st3) );
  ffd_async_274 wf1_cw3 ( .clk(clk), .reset(n33), .en(1'b1), .d(wf1_st2), .q(
        wf1_st3) );
  ffd_async_273 s3_cw4 ( .clk(clk), .reset(n33), .en(1'b1), .d(s3_st3), .q(
        s3_st4) );
  ffd_async_272 wf1_cw4 ( .clk(clk), .reset(n33), .en(1'b1), .d(wf1_st3), .q(
        wf1_st4) );
  NOR2_X2 U32 ( .A1(n30), .A2(n15), .ZN(inp2[15]) );
  NOR4_X2 U45 ( .A1(ir_st1[27]), .A2(ir_st1[28]), .A3(ir_st1[26]), .A4(n31), 
        .ZN(n30) );
  NOR2_X1 U3 ( .A1(n26), .A2(n25), .ZN(rd2[0]) );
  NOR2_X1 U4 ( .A1(n26), .A2(n19), .ZN(rd2[3]) );
  INV_X1 U5 ( .A(n30), .ZN(n14) );
  NOR2_X1 U6 ( .A1(n26), .A2(n17), .ZN(rd2[4]) );
  NOR2_X1 U7 ( .A1(n26), .A2(n21), .ZN(rd2[2]) );
  NOR2_X1 U8 ( .A1(n26), .A2(n23), .ZN(rd2[1]) );
  INV_X1 U9 ( .A(n16), .ZN(n26) );
  OAI22_X1 U10 ( .A1(n14), .A2(n24), .B1(n16), .B2(n25), .ZN(rd[0]) );
  OAI22_X1 U11 ( .A1(n14), .A2(n22), .B1(n16), .B2(n23), .ZN(rd[1]) );
  OAI22_X1 U12 ( .A1(n14), .A2(n20), .B1(n16), .B2(n21), .ZN(rd[2]) );
  OAI22_X1 U13 ( .A1(n14), .A2(n18), .B1(n16), .B2(n19), .ZN(rd[3]) );
  OAI22_X1 U14 ( .A1(n14), .A2(n15), .B1(n16), .B2(n17), .ZN(rd[4]) );
  NOR2_X1 U15 ( .A1(n30), .A2(n24), .ZN(inp2[11]) );
  NOR2_X1 U16 ( .A1(n30), .A2(n22), .ZN(inp2[12]) );
  NOR2_X1 U17 ( .A1(n30), .A2(n20), .ZN(inp2[13]) );
  NOR2_X1 U18 ( .A1(n30), .A2(n18), .ZN(inp2[14]) );
  BUF_X2 U19 ( .A(rst), .Z(n32) );
  BUF_X2 U20 ( .A(rst), .Z(n33) );
  OR3_X1 U21 ( .A1(ir_st1[29]), .A2(ir_st1[31]), .A3(ir_st1[30]), .ZN(n31) );
  NAND2_X1 U22 ( .A1(n14), .A2(n27), .ZN(n16) );
  NAND4_X1 U23 ( .A1(ir_st1[29]), .A2(ir_st1[27]), .A3(ir_st1[31]), .A4(n28), 
        .ZN(n27) );
  NOR3_X1 U24 ( .A1(n29), .A2(ir_st1[30]), .A3(ir_st1[28]), .ZN(n28) );
  INV_X1 U25 ( .A(ir_st1[26]), .ZN(n29) );
  INV_X1 U26 ( .A(ir_st1[18]), .ZN(n21) );
  INV_X1 U27 ( .A(ir_st1[20]), .ZN(n17) );
  INV_X1 U28 ( .A(ir_st1[17]), .ZN(n23) );
  INV_X1 U29 ( .A(ir_st1[19]), .ZN(n19) );
  INV_X1 U30 ( .A(ir_st1[16]), .ZN(n25) );
  INV_X1 U31 ( .A(ir_st1[11]), .ZN(n24) );
  INV_X1 U33 ( .A(ir_st1[12]), .ZN(n22) );
  INV_X1 U34 ( .A(ir_st1[13]), .ZN(n20) );
  INV_X1 U35 ( .A(ir_st1[14]), .ZN(n18) );
  INV_X1 U36 ( .A(ir_st1[15]), .ZN(n15) );
  AND2_X1 U37 ( .A1(ir_st1[0]), .A2(n14), .ZN(inp2[0]) );
  AND2_X1 U38 ( .A1(ir_st1[1]), .A2(n14), .ZN(inp2[1]) );
  AND2_X1 U39 ( .A1(ir_st1[2]), .A2(n14), .ZN(inp2[2]) );
  AND2_X1 U40 ( .A1(ir_st1[3]), .A2(n14), .ZN(inp2[3]) );
  AND2_X1 U41 ( .A1(ir_st1[4]), .A2(n14), .ZN(inp2[4]) );
  AND2_X1 U42 ( .A1(ir_st1[5]), .A2(n14), .ZN(inp2[5]) );
  AND2_X1 U43 ( .A1(ir_st1[6]), .A2(n14), .ZN(inp2[6]) );
  AND2_X1 U44 ( .A1(ir_st1[7]), .A2(n14), .ZN(inp2[7]) );
  AND2_X1 U46 ( .A1(ir_st1[8]), .A2(n14), .ZN(inp2[8]) );
  AND2_X1 U47 ( .A1(ir_st1[9]), .A2(n14), .ZN(inp2[9]) );
  AND2_X1 U48 ( .A1(ir_st1[10]), .A2(n14), .ZN(inp2[10]) );
endmodule


module CU_HW_OP_CODE_SIZE6_IR_SIZE32_FUNC_SIZE11_CW_SIZE18 ( Clk, Rst, IR_IN, 
        EN0, EN1, RF1, RF2, EN2, S1, S2, ALU1, ALU2, ALU3, ALU4, EQ_COND, 
        JUMP_EN, EN3, DEN, RW, S3, WF1 );
  input [31:0] IR_IN;
  input Clk, Rst;
  output EN0, EN1, RF1, RF2, EN2, S1, S2, ALU1, ALU2, ALU3, ALU4, EQ_COND,
         JUMP_EN, EN3, DEN, RW, S3, WF1;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26, N814, n1,
         n43, n44, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125;
  wire   [17:0] CW;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];

  DFF_X1 EN0_reg ( .D(CW[17]), .CK(N814), .Q(EN0), .QN(n1) );
  DFF_X1 EN1_reg ( .D(CW[4]), .CK(N814), .Q(EN1) );
  DFF_X1 RF1_reg ( .D(CW[15]), .CK(N814), .Q(RF1) );
  DFF_X1 RF2_reg ( .D(CW[14]), .CK(N814), .Q(RF2) );
  DFF_X1 EN2_reg ( .D(CW[4]), .CK(N814), .Q(EN2) );
  DFF_X1 S1_reg ( .D(CW[12]), .CK(N814), .Q(S1) );
  DFF_X1 S2_reg ( .D(CW[11]), .CK(N814), .Q(S2) );
  DFF_X1 ALU1_reg ( .D(CW[10]), .CK(N814), .Q(ALU1) );
  DFF_X1 ALU2_reg ( .D(CW[9]), .CK(N814), .Q(ALU2) );
  DFF_X1 ALU3_reg ( .D(CW[8]), .CK(N814), .Q(ALU3) );
  DFF_X1 ALU4_reg ( .D(CW[7]), .CK(N814), .Q(ALU4) );
  DFF_X1 EQ_COND_reg ( .D(CW[6]), .CK(N814), .Q(EQ_COND) );
  DFF_X1 JUMP_EN_reg ( .D(CW[5]), .CK(N814), .Q(JUMP_EN) );
  DFF_X1 EN3_reg ( .D(CW[4]), .CK(N814), .Q(EN3) );
  DFF_X1 DEN_reg ( .D(CW[3]), .CK(N814), .Q(DEN) );
  DFF_X1 RW_reg ( .D(CW[2]), .CK(N814), .Q(RW) );
  DFF_X1 S3_reg ( .D(CW[1]), .CK(N814), .Q(S3) );
  DFF_X1 WF1_reg ( .D(CW[0]), .CK(N814), .Q(WF1) );
  NAND3_X1 U91 ( .A1(n71), .A2(n79), .A3(n80), .ZN(CW[15]) );
  NAND3_X1 U92 ( .A1(n63), .A2(n49), .A3(n83), .ZN(n82) );
  NAND3_X1 U93 ( .A1(n71), .A2(n79), .A3(n84), .ZN(CW[12]) );
  NAND3_X1 U94 ( .A1(IR_IN_27), .A2(n92), .A3(n93), .ZN(n86) );
  NAND3_X1 U95 ( .A1(n89), .A2(IR_IN_30), .A3(n66), .ZN(n85) );
  NAND3_X1 U96 ( .A1(n65), .A2(n92), .A3(IR_IN_30), .ZN(n47) );
  NAND3_X1 U97 ( .A1(IR_IN_29), .A2(n104), .A3(n93), .ZN(n101) );
  NAND3_X1 U98 ( .A1(IR_IN_26), .A2(n90), .A3(n106), .ZN(n108) );
  NAND3_X1 U99 ( .A1(n116), .A2(n117), .A3(n112), .ZN(n110) );
  NAND3_X1 U100 ( .A1(IR_IN[2]), .A2(IR_IN[1]), .A3(n118), .ZN(n49) );
  NAND3_X1 U101 ( .A1(n120), .A2(n121), .A3(n122), .ZN(n115) );
  INV_X1 U3 ( .A(n71), .ZN(CW[1]) );
  AOI21_X1 U4 ( .B1(Rst), .B2(n78), .A(CW[6]), .ZN(n80) );
  NAND2_X1 U5 ( .A1(Rst), .A2(n74), .ZN(n71) );
  NOR2_X1 U6 ( .A1(n70), .A2(n125), .ZN(CW[4]) );
  NAND2_X1 U7 ( .A1(n70), .A2(Rst), .ZN(CW[17]) );
  OAI21_X1 U8 ( .B1(n73), .B2(n52), .A(Rst), .ZN(n84) );
  INV_X1 U9 ( .A(n79), .ZN(CW[3]) );
  AND2_X1 U10 ( .A1(n77), .A2(Rst), .ZN(CW[6]) );
  NAND2_X1 U11 ( .A1(n94), .A2(n71), .ZN(CW[0]) );
  INV_X1 U12 ( .A(n94), .ZN(CW[2]) );
  NOR4_X1 U13 ( .A1(n72), .A2(n73), .A3(n74), .A4(n75), .ZN(n70) );
  OR4_X1 U14 ( .A1(n76), .A2(n77), .A3(n78), .A4(n52), .ZN(n75) );
  AOI21_X1 U15 ( .B1(Rst), .B2(n72), .A(CW[2]), .ZN(n79) );
  NOR2_X1 U16 ( .A1(n54), .A2(n125), .ZN(CW[8]) );
  NOR3_X1 U17 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n54) );
  OR3_X1 U18 ( .A1(n58), .A2(n52), .A3(n51), .ZN(n55) );
  NOR2_X1 U19 ( .A1(n81), .A2(n125), .ZN(CW[14]) );
  NOR3_X1 U20 ( .A1(n82), .A2(n72), .A3(n56), .ZN(n81) );
  OAI21_X1 U21 ( .B1(n105), .B2(n90), .A(n46), .ZN(n57) );
  AOI211_X1 U22 ( .C1(n91), .C2(n89), .A(n67), .B(n106), .ZN(n105) );
  NAND4_X1 U23 ( .A1(n63), .A2(n49), .A3(n83), .A4(n99), .ZN(n74) );
  NOR2_X1 U24 ( .A1(n56), .A2(n88), .ZN(n99) );
  NOR2_X1 U25 ( .A1(n51), .A2(n106), .ZN(n98) );
  OAI21_X1 U26 ( .B1(n125), .B2(n86), .A(n80), .ZN(CW[5]) );
  INV_X1 U27 ( .A(n85), .ZN(n52) );
  NAND2_X1 U28 ( .A1(n114), .A2(n112), .ZN(n83) );
  NAND2_X1 U29 ( .A1(n76), .A2(Rst), .ZN(n94) );
  INV_X1 U30 ( .A(n115), .ZN(n113) );
  INV_X1 U31 ( .A(n63), .ZN(n58) );
  INV_X1 U32 ( .A(n86), .ZN(n73) );
  AND3_X1 U33 ( .A1(n89), .A2(n90), .A3(n91), .ZN(n78) );
  AND3_X1 U34 ( .A1(n89), .A2(n90), .A3(n66), .ZN(n77) );
  INV_X1 U35 ( .A(n93), .ZN(n123) );
  INV_X1 U36 ( .A(n91), .ZN(n124) );
  OR2_X1 U37 ( .A1(n66), .A2(n91), .ZN(n92) );
  INV_X1 U38 ( .A(n64), .ZN(n61) );
  AOI21_X1 U39 ( .B1(n65), .B2(n66), .A(n67), .ZN(n64) );
  INV_X1 U40 ( .A(n87), .ZN(CW[11]) );
  AOI211_X1 U41 ( .C1(n88), .C2(Rst), .A(CW[3]), .B(CW[5]), .ZN(n87) );
  INV_X1 U42 ( .A(Rst), .ZN(n125) );
  NOR4_X1 U43 ( .A1(n104), .A2(n107), .A3(IR_IN_27), .A4(IR_IN_31), .ZN(n67)
         );
  INV_X1 U44 ( .A(IR_IN_29), .ZN(n107) );
  NOR3_X1 U45 ( .A1(IR_IN_27), .A2(IR_IN_31), .A3(n103), .ZN(n89) );
  OAI221_X1 U46 ( .B1(n110), .B2(n111), .C1(n112), .C2(n53), .A(n48), .ZN(n56)
         );
  NAND2_X1 U47 ( .A1(IR_IN[2]), .A2(n113), .ZN(n111) );
  INV_X1 U48 ( .A(IR_IN[1]), .ZN(n116) );
  NOR3_X1 U49 ( .A1(n115), .A2(IR_IN[1]), .A3(n117), .ZN(n114) );
  NOR3_X1 U50 ( .A1(n115), .A2(IR_IN[5]), .A3(IR_IN[3]), .ZN(n118) );
  NOR3_X1 U51 ( .A1(IR_IN_30), .A2(IR_IN_31), .A3(IR_IN_28), .ZN(n93) );
  NAND4_X1 U52 ( .A1(IR_IN_29), .A2(IR_IN_27), .A3(n109), .A4(n104), .ZN(n46)
         );
  NOR2_X1 U53 ( .A1(IR_IN_31), .A2(IR_IN_30), .ZN(n109) );
  NOR2_X1 U54 ( .A1(IR_IN[3]), .A2(IR_IN[0]), .ZN(n112) );
  NOR3_X1 U55 ( .A1(n102), .A2(IR_IN_30), .A3(IR_IN_28), .ZN(n95) );
  NOR2_X1 U56 ( .A1(n104), .A2(IR_IN_29), .ZN(n66) );
  OAI21_X1 U57 ( .B1(IR_IN_28), .B2(n46), .A(n108), .ZN(n51) );
  NAND4_X1 U58 ( .A1(IR_IN[5]), .A2(IR_IN[1]), .A3(n113), .A4(n112), .ZN(n48)
         );
  NOR2_X1 U59 ( .A1(IR_IN[7]), .A2(IR_IN[6]), .ZN(n120) );
  NOR3_X1 U60 ( .A1(IR_IN[8]), .A2(IR_IN_27), .A3(IR_IN[9]), .ZN(n121) );
  NOR4_X1 U61 ( .A1(IR_IN[4]), .A2(IR_IN[10]), .A3(n123), .A4(n124), .ZN(n122)
         );
  NOR3_X1 U62 ( .A1(n102), .A2(IR_IN_31), .A3(n103), .ZN(n65) );
  NOR2_X1 U63 ( .A1(IR_IN_26), .A2(IR_IN_29), .ZN(n91) );
  NAND4_X1 U64 ( .A1(IR_IN[3]), .A2(IR_IN[0]), .A3(n114), .A4(n119), .ZN(n63)
         );
  INV_X1 U65 ( .A(IR_IN[2]), .ZN(n119) );
  NAND4_X1 U66 ( .A1(n98), .A2(n100), .A3(n101), .A4(n47), .ZN(n88) );
  INV_X1 U67 ( .A(n57), .ZN(n100) );
  NAND2_X1 U68 ( .A1(n114), .A2(IR_IN[2]), .ZN(n53) );
  INV_X1 U69 ( .A(IR_IN_26), .ZN(n104) );
  AOI21_X1 U70 ( .B1(n59), .B2(n60), .A(n125), .ZN(CW[7]) );
  INV_X1 U71 ( .A(n68), .ZN(n59) );
  AOI221_X1 U72 ( .B1(IR_IN_30), .B2(n61), .C1(n62), .C2(IR_IN[3]), .A(n58), 
        .ZN(n60) );
  OAI222_X1 U73 ( .A1(n46), .A2(IR_IN_28), .B1(n49), .B2(n69), .C1(n48), .C2(
        IR_IN[2]), .ZN(n68) );
  INV_X1 U74 ( .A(IR_IN_30), .ZN(n90) );
  NOR2_X1 U75 ( .A1(IR_IN[0]), .A2(n53), .ZN(n62) );
  AOI21_X1 U76 ( .B1(n43), .B2(n44), .A(n125), .ZN(CW[9]) );
  AND4_X1 U77 ( .A1(n46), .A2(n47), .A3(n48), .A4(n49), .ZN(n44) );
  AOI211_X1 U78 ( .C1(n50), .C2(IR_IN[0]), .A(n51), .B(n52), .ZN(n43) );
  NOR2_X1 U79 ( .A1(IR_IN[3]), .A2(n53), .ZN(n50) );
  AND2_X1 U80 ( .A1(n89), .A2(IR_IN_29), .ZN(n106) );
  INV_X1 U81 ( .A(IR_IN_27), .ZN(n102) );
  AND4_X1 U82 ( .A1(IR_IN_26), .A2(IR_IN_29), .A3(IR_IN_31), .A4(n95), .ZN(n72) );
  INV_X1 U83 ( .A(IR_IN_28), .ZN(n103) );
  AND3_X1 U84 ( .A1(IR_IN_31), .A2(n66), .A3(n95), .ZN(n76) );
  INV_X1 U85 ( .A(IR_IN[5]), .ZN(n117) );
  AND2_X1 U86 ( .A1(n96), .A2(Rst), .ZN(CW[10]) );
  OAI211_X1 U87 ( .C1(n48), .C2(IR_IN[2]), .A(n97), .B(n98), .ZN(n96) );
  AND2_X1 U88 ( .A1(n85), .A2(n53), .ZN(n97) );
  INV_X1 U89 ( .A(IR_IN[0]), .ZN(n69) );
  INV_X1 U90 ( .A(Clk), .ZN(N814) );
endmodule


module DLX_IR_SIZE32_PC_SIZE32 ( CLK, RST, IRAM_ADDRESS, IRAM_ISSUE, 
        IRAM_READY, IRAM_DATA, DRAM_ADDRESS, DRAM_READNOTWRITE, DRAM_ISSUE, 
        DRAM_DATA_in, DRAM_READY, DRAM_DATA_out );
  output [31:0] IRAM_ADDRESS;
  input [31:0] IRAM_DATA;
  output [31:0] DRAM_ADDRESS;
  input [31:0] DRAM_DATA_in;
  output [31:0] DRAM_DATA_out;
  input CLK, RST, IRAM_READY, DRAM_READY;
  output IRAM_ISSUE, DRAM_READNOTWRITE, DRAM_ISSUE;
  wire   EN0_int, EN1_int, RF1_int, RF2_int, EN2_int, S1_int, S2_int, ALU1_int,
         ALU2_int, ALU3_int, ALU4_int, EQ_COND_int, JUMP_EN_int, EN3_int,
         DEN_int, RW_int, S3_int, WF1_int, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382;
  wire   [31:0] IR;
  wire   [31:0] pc_in_i;
  wire   [31:0] pc_out_i;

  DFFR_X1 \IR_reg[0]  ( .D(n257), .CK(CLK), .RN(n376), .Q(IR[0]), .QN(n161) );
  DFFR_X1 \IR_reg[1]  ( .D(n256), .CK(CLK), .RN(n382), .Q(IR[1]), .QN(n160) );
  DFFR_X1 \IR_reg[2]  ( .D(n255), .CK(CLK), .RN(n382), .Q(IR[2]), .QN(n159) );
  DFFR_X1 \IR_reg[3]  ( .D(n254), .CK(CLK), .RN(n382), .Q(IR[3]), .QN(n158) );
  DFFR_X1 \IR_reg[4]  ( .D(n253), .CK(CLK), .RN(n382), .Q(IR[4]), .QN(n157) );
  DFFR_X1 \IR_reg[5]  ( .D(n252), .CK(CLK), .RN(n382), .Q(IR[5]), .QN(n156) );
  DFFR_X1 \IR_reg[6]  ( .D(n251), .CK(CLK), .RN(n381), .Q(IR[6]), .QN(n155) );
  DFFR_X1 \IR_reg[7]  ( .D(n250), .CK(CLK), .RN(n381), .Q(IR[7]), .QN(n154) );
  DFFR_X1 \IR_reg[8]  ( .D(n249), .CK(CLK), .RN(n381), .Q(IR[8]), .QN(n153) );
  DFFR_X1 \IR_reg[9]  ( .D(n248), .CK(CLK), .RN(n381), .Q(IR[9]), .QN(n152) );
  DFFR_X1 \IR_reg[10]  ( .D(n247), .CK(CLK), .RN(n381), .Q(IR[10]), .QN(n151)
         );
  DFFR_X1 \IR_reg[11]  ( .D(n246), .CK(CLK), .RN(n381), .Q(IR[11]), .QN(n150)
         );
  DFFR_X1 \IR_reg[12]  ( .D(n245), .CK(CLK), .RN(n381), .Q(IR[12]), .QN(n149)
         );
  DFFR_X1 \IR_reg[13]  ( .D(n244), .CK(CLK), .RN(n381), .Q(IR[13]), .QN(n148)
         );
  DFFR_X1 \IR_reg[14]  ( .D(n243), .CK(CLK), .RN(n381), .Q(IR[14]), .QN(n147)
         );
  DFFR_X1 \IR_reg[15]  ( .D(n242), .CK(CLK), .RN(n381), .Q(IR[15]), .QN(n146)
         );
  DFFR_X1 \IR_reg[16]  ( .D(n241), .CK(CLK), .RN(n381), .Q(IR[16]), .QN(n145)
         );
  DFFR_X1 \IR_reg[17]  ( .D(n240), .CK(CLK), .RN(n381), .Q(IR[17]), .QN(n144)
         );
  DFFR_X1 \IR_reg[18]  ( .D(n239), .CK(CLK), .RN(n381), .Q(IR[18]), .QN(n143)
         );
  DFFR_X1 \IR_reg[19]  ( .D(n238), .CK(CLK), .RN(n381), .Q(IR[19]), .QN(n142)
         );
  DFFR_X1 \IR_reg[20]  ( .D(n237), .CK(CLK), .RN(n381), .Q(IR[20]), .QN(n141)
         );
  DFFR_X1 \IR_reg[21]  ( .D(n236), .CK(CLK), .RN(n381), .Q(IR[21]), .QN(n140)
         );
  DFFR_X1 \IR_reg[22]  ( .D(n235), .CK(CLK), .RN(n380), .Q(IR[22]), .QN(n139)
         );
  DFFR_X1 \IR_reg[23]  ( .D(n234), .CK(CLK), .RN(n380), .Q(IR[23]), .QN(n138)
         );
  DFFR_X1 \IR_reg[24]  ( .D(n233), .CK(CLK), .RN(n380), .Q(IR[24]), .QN(n137)
         );
  DFFR_X1 \IR_reg[25]  ( .D(n232), .CK(CLK), .RN(n380), .Q(IR[25]), .QN(n136)
         );
  DFFR_X1 \IR_reg[26]  ( .D(n231), .CK(CLK), .RN(n380), .Q(IR[26]), .QN(n135)
         );
  DFFR_X1 \IR_reg[27]  ( .D(n230), .CK(CLK), .RN(n380), .Q(IR[27]), .QN(n134)
         );
  DFFR_X1 \IR_reg[28]  ( .D(n229), .CK(CLK), .RN(n380), .Q(IR[28]), .QN(n133)
         );
  DFFR_X1 \IR_reg[29]  ( .D(n228), .CK(CLK), .RN(n380), .Q(IR[29]), .QN(n132)
         );
  DFFR_X1 \IR_reg[30]  ( .D(n227), .CK(CLK), .RN(n380), .Q(IR[30]), .QN(n131)
         );
  DFFR_X1 \IR_reg[31]  ( .D(n226), .CK(CLK), .RN(n380), .Q(IR[31]), .QN(n130)
         );
  DFFR_X1 \pc_in_i_reg[0]  ( .D(n225), .CK(CLK), .RN(n380), .Q(pc_in_i[0]), 
        .QN(n66) );
  DFFR_X1 \IRAM_ADDRESS_reg[0]  ( .D(n224), .CK(CLK), .RN(n380), .Q(
        IRAM_ADDRESS[0]), .QN(n129) );
  DFFR_X1 \pc_in_i_reg[1]  ( .D(n223), .CK(CLK), .RN(n380), .Q(pc_in_i[1]), 
        .QN(n67) );
  DFFR_X1 \IRAM_ADDRESS_reg[1]  ( .D(n222), .CK(CLK), .RN(n376), .Q(
        IRAM_ADDRESS[1]), .QN(n128) );
  DFFR_X1 \pc_in_i_reg[2]  ( .D(n221), .CK(CLK), .RN(n380), .Q(pc_in_i[2]), 
        .QN(n68) );
  DFFR_X1 \IRAM_ADDRESS_reg[2]  ( .D(n220), .CK(CLK), .RN(n380), .Q(
        IRAM_ADDRESS[2]), .QN(n127) );
  DFFR_X1 \pc_in_i_reg[3]  ( .D(n219), .CK(CLK), .RN(n379), .Q(pc_in_i[3]), 
        .QN(n69) );
  DFFR_X1 \IRAM_ADDRESS_reg[3]  ( .D(n218), .CK(CLK), .RN(n379), .Q(
        IRAM_ADDRESS[3]), .QN(n126) );
  DFFR_X1 \pc_in_i_reg[4]  ( .D(n217), .CK(CLK), .RN(n379), .Q(pc_in_i[4]), 
        .QN(n70) );
  DFFR_X1 \IRAM_ADDRESS_reg[4]  ( .D(n216), .CK(CLK), .RN(n379), .Q(
        IRAM_ADDRESS[4]), .QN(n125) );
  DFFR_X1 \pc_in_i_reg[5]  ( .D(n215), .CK(CLK), .RN(n379), .Q(pc_in_i[5]), 
        .QN(n71) );
  DFFR_X1 \IRAM_ADDRESS_reg[5]  ( .D(n214), .CK(CLK), .RN(n379), .Q(
        IRAM_ADDRESS[5]), .QN(n124) );
  DFFR_X1 \pc_in_i_reg[6]  ( .D(n213), .CK(CLK), .RN(n379), .Q(pc_in_i[6]), 
        .QN(n72) );
  DFFR_X1 \IRAM_ADDRESS_reg[6]  ( .D(n212), .CK(CLK), .RN(n379), .Q(
        IRAM_ADDRESS[6]), .QN(n123) );
  DFFR_X1 \pc_in_i_reg[7]  ( .D(n211), .CK(CLK), .RN(n379), .Q(pc_in_i[7]), 
        .QN(n73) );
  DFFR_X1 \IRAM_ADDRESS_reg[7]  ( .D(n210), .CK(CLK), .RN(n379), .Q(
        IRAM_ADDRESS[7]), .QN(n122) );
  DFFR_X1 \pc_in_i_reg[8]  ( .D(n209), .CK(CLK), .RN(n379), .Q(pc_in_i[8]), 
        .QN(n74) );
  DFFR_X1 \IRAM_ADDRESS_reg[8]  ( .D(n208), .CK(CLK), .RN(n379), .Q(
        IRAM_ADDRESS[8]), .QN(n121) );
  DFFR_X1 \pc_in_i_reg[9]  ( .D(n207), .CK(CLK), .RN(n379), .Q(pc_in_i[9]), 
        .QN(n75) );
  DFFR_X1 \IRAM_ADDRESS_reg[9]  ( .D(n206), .CK(CLK), .RN(n379), .Q(
        IRAM_ADDRESS[9]), .QN(n120) );
  DFFR_X1 \pc_in_i_reg[10]  ( .D(n205), .CK(CLK), .RN(n379), .Q(pc_in_i[10]), 
        .QN(n76) );
  DFFR_X1 \IRAM_ADDRESS_reg[10]  ( .D(n204), .CK(CLK), .RN(n378), .Q(
        IRAM_ADDRESS[10]), .QN(n119) );
  DFFR_X1 \pc_in_i_reg[11]  ( .D(n203), .CK(CLK), .RN(n378), .Q(pc_in_i[11]), 
        .QN(n77) );
  DFFR_X1 \IRAM_ADDRESS_reg[11]  ( .D(n202), .CK(CLK), .RN(n378), .Q(
        IRAM_ADDRESS[11]), .QN(n118) );
  DFFR_X1 \pc_in_i_reg[12]  ( .D(n201), .CK(CLK), .RN(n378), .Q(pc_in_i[12]), 
        .QN(n78) );
  DFFR_X1 \IRAM_ADDRESS_reg[12]  ( .D(n200), .CK(CLK), .RN(n378), .Q(
        IRAM_ADDRESS[12]), .QN(n117) );
  DFFR_X1 \pc_in_i_reg[13]  ( .D(n199), .CK(CLK), .RN(n378), .Q(pc_in_i[13]), 
        .QN(n79) );
  DFFR_X1 \IRAM_ADDRESS_reg[13]  ( .D(n198), .CK(CLK), .RN(n378), .Q(
        IRAM_ADDRESS[13]), .QN(n116) );
  DFFR_X1 \pc_in_i_reg[14]  ( .D(n197), .CK(CLK), .RN(n378), .Q(pc_in_i[14]), 
        .QN(n80) );
  DFFR_X1 \IRAM_ADDRESS_reg[14]  ( .D(n196), .CK(CLK), .RN(n378), .Q(
        IRAM_ADDRESS[14]), .QN(n115) );
  DFFR_X1 \pc_in_i_reg[15]  ( .D(n195), .CK(CLK), .RN(n378), .Q(pc_in_i[15]), 
        .QN(n81) );
  DFFR_X1 \IRAM_ADDRESS_reg[15]  ( .D(n194), .CK(CLK), .RN(n378), .Q(
        IRAM_ADDRESS[15]), .QN(n114) );
  DFFR_X1 \pc_in_i_reg[16]  ( .D(n193), .CK(CLK), .RN(n378), .Q(pc_in_i[16]), 
        .QN(n82) );
  DFFR_X1 \IRAM_ADDRESS_reg[16]  ( .D(n192), .CK(CLK), .RN(n378), .Q(
        IRAM_ADDRESS[16]), .QN(n113) );
  DFFR_X1 \pc_in_i_reg[17]  ( .D(n191), .CK(CLK), .RN(n378), .Q(pc_in_i[17]), 
        .QN(n83) );
  DFFR_X1 \IRAM_ADDRESS_reg[17]  ( .D(n190), .CK(CLK), .RN(n378), .Q(
        IRAM_ADDRESS[17]), .QN(n112) );
  DFFR_X1 \pc_in_i_reg[18]  ( .D(n189), .CK(CLK), .RN(n378), .Q(pc_in_i[18]), 
        .QN(n84) );
  DFFR_X1 \IRAM_ADDRESS_reg[18]  ( .D(n188), .CK(CLK), .RN(n377), .Q(
        IRAM_ADDRESS[18]), .QN(n111) );
  DFFR_X1 \pc_in_i_reg[19]  ( .D(n187), .CK(CLK), .RN(n377), .Q(pc_in_i[19]), 
        .QN(n85) );
  DFFR_X1 \IRAM_ADDRESS_reg[19]  ( .D(n186), .CK(CLK), .RN(n377), .Q(
        IRAM_ADDRESS[19]), .QN(n110) );
  DFFR_X1 \pc_in_i_reg[20]  ( .D(n185), .CK(CLK), .RN(n377), .Q(pc_in_i[20]), 
        .QN(n86) );
  DFFR_X1 \IRAM_ADDRESS_reg[20]  ( .D(n184), .CK(CLK), .RN(n379), .Q(
        IRAM_ADDRESS[20]), .QN(n109) );
  DFFR_X1 \pc_in_i_reg[21]  ( .D(n183), .CK(CLK), .RN(n377), .Q(pc_in_i[21]), 
        .QN(n87) );
  DFFR_X1 \IRAM_ADDRESS_reg[21]  ( .D(n182), .CK(CLK), .RN(n377), .Q(
        IRAM_ADDRESS[21]), .QN(n108) );
  DFFR_X1 \pc_in_i_reg[22]  ( .D(n181), .CK(CLK), .RN(n377), .Q(pc_in_i[22]), 
        .QN(n88) );
  DFFR_X1 \IRAM_ADDRESS_reg[22]  ( .D(n180), .CK(CLK), .RN(n377), .Q(
        IRAM_ADDRESS[22]), .QN(n107) );
  DFFR_X1 \pc_in_i_reg[23]  ( .D(n179), .CK(CLK), .RN(n377), .Q(pc_in_i[23]), 
        .QN(n89) );
  DFFR_X1 \IRAM_ADDRESS_reg[23]  ( .D(n178), .CK(CLK), .RN(n377), .Q(
        IRAM_ADDRESS[23]), .QN(n106) );
  DFFR_X1 \pc_in_i_reg[24]  ( .D(n177), .CK(CLK), .RN(n377), .Q(pc_in_i[24]), 
        .QN(n90) );
  DFFR_X1 \IRAM_ADDRESS_reg[24]  ( .D(n176), .CK(CLK), .RN(n377), .Q(
        IRAM_ADDRESS[24]), .QN(n105) );
  DFFR_X1 \pc_in_i_reg[25]  ( .D(n175), .CK(CLK), .RN(n377), .Q(pc_in_i[25]), 
        .QN(n91) );
  DFFR_X1 \IRAM_ADDRESS_reg[25]  ( .D(n174), .CK(CLK), .RN(n377), .Q(
        IRAM_ADDRESS[25]), .QN(n104) );
  DFFR_X1 \pc_in_i_reg[26]  ( .D(n173), .CK(CLK), .RN(n377), .Q(pc_in_i[26]), 
        .QN(n92) );
  DFFR_X1 \IRAM_ADDRESS_reg[26]  ( .D(n172), .CK(CLK), .RN(n377), .Q(
        IRAM_ADDRESS[26]), .QN(n103) );
  DFFR_X1 \pc_in_i_reg[27]  ( .D(n171), .CK(CLK), .RN(n376), .Q(pc_in_i[27]), 
        .QN(n93) );
  DFFR_X1 \IRAM_ADDRESS_reg[27]  ( .D(n170), .CK(CLK), .RN(n376), .Q(
        IRAM_ADDRESS[27]), .QN(n102) );
  DFFR_X1 \pc_in_i_reg[28]  ( .D(n169), .CK(CLK), .RN(n376), .Q(pc_in_i[28]), 
        .QN(n94) );
  DFFR_X1 \IRAM_ADDRESS_reg[28]  ( .D(n168), .CK(CLK), .RN(n376), .Q(
        IRAM_ADDRESS[28]), .QN(n101) );
  DFFR_X1 \pc_in_i_reg[29]  ( .D(n167), .CK(CLK), .RN(n376), .Q(pc_in_i[29]), 
        .QN(n95) );
  DFFR_X1 \IRAM_ADDRESS_reg[29]  ( .D(n166), .CK(CLK), .RN(n376), .Q(
        IRAM_ADDRESS[29]), .QN(n100) );
  DFFR_X1 \pc_in_i_reg[30]  ( .D(n165), .CK(CLK), .RN(n376), .Q(pc_in_i[30]), 
        .QN(n96) );
  DFFR_X1 \IRAM_ADDRESS_reg[30]  ( .D(n164), .CK(CLK), .RN(n376), .Q(
        IRAM_ADDRESS[30]), .QN(n99) );
  DFFR_X1 \pc_in_i_reg[31]  ( .D(n163), .CK(CLK), .RN(n380), .Q(pc_in_i[31]), 
        .QN(n97) );
  DFFR_X1 \IRAM_ADDRESS_reg[31]  ( .D(n162), .CK(CLK), .RN(n376), .Q(
        IRAM_ADDRESS[31]), .QN(n98) );
  CU_HW_OP_CODE_SIZE6_IR_SIZE32_FUNC_SIZE11_CW_SIZE18 CU ( .Clk(CLK), .Rst(
        n376), .IR_IN(IR), .EN0(EN0_int), .EN1(EN1_int), .RF1(RF1_int), .RF2(
        RF2_int), .EN2(EN2_int), .S1(S1_int), .S2(S2_int), .ALU1(ALU1_int), 
        .ALU2(ALU2_int), .ALU3(ALU3_int), .ALU4(ALU4_int), .EQ_COND(
        EQ_COND_int), .JUMP_EN(JUMP_EN_int), .EN3(EN3_int), .DEN(DEN_int), 
        .RW(RW_int), .S3(S3_int), .WF1(WF1_int) );
  datapath dp ( .clk(CLK), .rst(n376), .en0(n358), .ir(IR), .pc_in(pc_in_i), 
        .en1(EN1_int), .rf1(RF1_int), .rf2(RF2_int), .en2(EN2_int), .s1(S1_int), .s2(S2_int), .alu1(ALU1_int), .alu2(ALU2_int), .alu3(ALU3_int), .alu4(
        ALU4_int), .eq_cond(EQ_COND_int), .jump_en(JUMP_EN_int), .en3(EN3_int), 
        .rw(RW_int), .den(DEN_int), .dram_data_in(DRAM_DATA_in), .dram_rw_en(
        DRAM_READNOTWRITE), .dram_enable(DRAM_ISSUE), .dram_data_out(
        DRAM_DATA_out), .dram_addr(DRAM_ADDRESS), .pc_out(pc_out_i), .s3(
        S3_int), .wf1(WF1_int) );
  INV_X1 U324 ( .A(n374), .ZN(n360) );
  INV_X1 U325 ( .A(n374), .ZN(n359) );
  INV_X1 U326 ( .A(n374), .ZN(n358) );
  BUF_X1 U327 ( .A(n375), .Z(n374) );
  BUF_X1 U328 ( .A(n375), .Z(n373) );
  BUF_X1 U329 ( .A(n371), .Z(n372) );
  BUF_X1 U330 ( .A(n375), .Z(n371) );
  BUF_X1 U331 ( .A(n368), .Z(n370) );
  BUF_X1 U332 ( .A(n375), .Z(n369) );
  BUF_X1 U333 ( .A(n375), .Z(n368) );
  BUF_X1 U334 ( .A(n375), .Z(n367) );
  BUF_X1 U335 ( .A(n367), .Z(n366) );
  BUF_X1 U336 ( .A(n369), .Z(n365) );
  BUF_X1 U337 ( .A(n368), .Z(n364) );
  BUF_X1 U338 ( .A(n372), .Z(n363) );
  BUF_X1 U339 ( .A(n365), .Z(n362) );
  BUF_X1 U340 ( .A(n367), .Z(n361) );
  INV_X1 U341 ( .A(n356), .ZN(n375) );
  OAI22_X1 U342 ( .A1(n373), .A2(n355), .B1(n98), .B2(n357), .ZN(n162) );
  OAI22_X1 U343 ( .A1(n373), .A2(n354), .B1(n99), .B2(n360), .ZN(n164) );
  OAI22_X1 U344 ( .A1(n371), .A2(n349), .B1(n104), .B2(n359), .ZN(n174) );
  OAI22_X1 U345 ( .A1(n369), .A2(n345), .B1(n108), .B2(n358), .ZN(n182) );
  OAI22_X1 U346 ( .A1(n372), .A2(n353), .B1(n100), .B2(n360), .ZN(n166) );
  OAI22_X1 U347 ( .A1(n372), .A2(n352), .B1(n101), .B2(n358), .ZN(n168) );
  OAI22_X1 U348 ( .A1(n372), .A2(n351), .B1(n102), .B2(n357), .ZN(n170) );
  OAI22_X1 U349 ( .A1(n371), .A2(n350), .B1(n103), .B2(n360), .ZN(n172) );
  OAI22_X1 U350 ( .A1(n370), .A2(n348), .B1(n105), .B2(n359), .ZN(n176) );
  OAI22_X1 U351 ( .A1(n370), .A2(n347), .B1(n106), .B2(n357), .ZN(n178) );
  OAI22_X1 U352 ( .A1(n370), .A2(n346), .B1(n107), .B2(n357), .ZN(n180) );
  OAI22_X1 U353 ( .A1(n369), .A2(n344), .B1(n109), .B2(n357), .ZN(n184) );
  OAI22_X1 U354 ( .A1(n368), .A2(n343), .B1(n110), .B2(n359), .ZN(n186) );
  OAI22_X1 U355 ( .A1(n368), .A2(n342), .B1(n111), .B2(EN0_int), .ZN(n188) );
  OAI22_X1 U356 ( .A1(n368), .A2(n341), .B1(n112), .B2(n357), .ZN(n190) );
  OAI22_X1 U357 ( .A1(n367), .A2(n340), .B1(n113), .B2(n357), .ZN(n192) );
  OAI22_X1 U358 ( .A1(n367), .A2(n339), .B1(n114), .B2(EN0_int), .ZN(n194) );
  OAI22_X1 U359 ( .A1(n366), .A2(n338), .B1(n115), .B2(n359), .ZN(n196) );
  OAI22_X1 U360 ( .A1(n366), .A2(n337), .B1(n116), .B2(n360), .ZN(n198) );
  OAI22_X1 U361 ( .A1(n365), .A2(n335), .B1(n118), .B2(n357), .ZN(n202) );
  OAI22_X1 U362 ( .A1(n365), .A2(n334), .B1(n119), .B2(n358), .ZN(n204) );
  OAI22_X1 U363 ( .A1(n364), .A2(n333), .B1(n120), .B2(n357), .ZN(n206) );
  OAI22_X1 U364 ( .A1(n364), .A2(n332), .B1(n121), .B2(n357), .ZN(n208) );
  OAI22_X1 U365 ( .A1(n364), .A2(n331), .B1(n122), .B2(n357), .ZN(n210) );
  OAI22_X1 U366 ( .A1(n363), .A2(n330), .B1(n123), .B2(n357), .ZN(n212) );
  OAI22_X1 U367 ( .A1(n363), .A2(n329), .B1(n124), .B2(n357), .ZN(n214) );
  OAI22_X1 U368 ( .A1(n362), .A2(n327), .B1(n126), .B2(n357), .ZN(n218) );
  OAI22_X1 U369 ( .A1(n362), .A2(n326), .B1(n127), .B2(n357), .ZN(n220) );
  OAI22_X1 U370 ( .A1(n366), .A2(n336), .B1(n117), .B2(n360), .ZN(n200) );
  OAI22_X1 U371 ( .A1(n362), .A2(n328), .B1(n125), .B2(n359), .ZN(n216) );
  OAI22_X1 U372 ( .A1(n361), .A2(n325), .B1(n128), .B2(n357), .ZN(n222) );
  OAI22_X1 U373 ( .A1(n361), .A2(n324), .B1(n129), .B2(n358), .ZN(n224) );
  OAI22_X1 U374 ( .A1(n371), .A2(n349), .B1(n360), .B2(n91), .ZN(n175) );
  OAI22_X1 U375 ( .A1(n370), .A2(n348), .B1(n360), .B2(n90), .ZN(n177) );
  OAI22_X1 U376 ( .A1(n370), .A2(n347), .B1(n360), .B2(n89), .ZN(n179) );
  OAI22_X1 U377 ( .A1(n369), .A2(n346), .B1(n360), .B2(n88), .ZN(n181) );
  OAI22_X1 U378 ( .A1(n369), .A2(n345), .B1(n360), .B2(n87), .ZN(n183) );
  OAI22_X1 U379 ( .A1(n369), .A2(n344), .B1(n360), .B2(n86), .ZN(n185) );
  OAI22_X1 U380 ( .A1(n368), .A2(n343), .B1(n360), .B2(n85), .ZN(n187) );
  OAI22_X1 U381 ( .A1(n368), .A2(n342), .B1(n360), .B2(n84), .ZN(n189) );
  OAI22_X1 U382 ( .A1(n367), .A2(n341), .B1(n360), .B2(n83), .ZN(n191) );
  OAI22_X1 U383 ( .A1(n367), .A2(n340), .B1(n359), .B2(n82), .ZN(n193) );
  OAI22_X1 U384 ( .A1(n367), .A2(n339), .B1(n360), .B2(n81), .ZN(n195) );
  OAI22_X1 U385 ( .A1(n366), .A2(n338), .B1(n360), .B2(n80), .ZN(n197) );
  OAI22_X1 U386 ( .A1(n366), .A2(n337), .B1(n360), .B2(n79), .ZN(n199) );
  OAI22_X1 U387 ( .A1(n365), .A2(n336), .B1(n360), .B2(n78), .ZN(n201) );
  OAI22_X1 U388 ( .A1(n365), .A2(n335), .B1(n359), .B2(n77), .ZN(n203) );
  OAI22_X1 U389 ( .A1(n365), .A2(n334), .B1(n359), .B2(n76), .ZN(n205) );
  OAI22_X1 U390 ( .A1(n364), .A2(n333), .B1(n359), .B2(n75), .ZN(n207) );
  OAI22_X1 U391 ( .A1(n364), .A2(n332), .B1(n359), .B2(n74), .ZN(n209) );
  OAI22_X1 U392 ( .A1(n363), .A2(n331), .B1(n359), .B2(n73), .ZN(n211) );
  OAI22_X1 U393 ( .A1(n363), .A2(n330), .B1(n359), .B2(n72), .ZN(n213) );
  OAI22_X1 U394 ( .A1(n363), .A2(n329), .B1(n359), .B2(n71), .ZN(n215) );
  OAI22_X1 U395 ( .A1(n362), .A2(n328), .B1(n359), .B2(n70), .ZN(n217) );
  OAI22_X1 U396 ( .A1(n362), .A2(n327), .B1(n359), .B2(n69), .ZN(n219) );
  OAI22_X1 U397 ( .A1(n361), .A2(n326), .B1(n359), .B2(n68), .ZN(n221) );
  OAI22_X1 U398 ( .A1(n361), .A2(n325), .B1(n359), .B2(n67), .ZN(n223) );
  OAI22_X1 U399 ( .A1(n361), .A2(n324), .B1(n359), .B2(n66), .ZN(n225) );
  OAI22_X1 U400 ( .A1(n373), .A2(n355), .B1(n356), .B2(n97), .ZN(n163) );
  OAI22_X1 U401 ( .A1(n373), .A2(n354), .B1(n357), .B2(n96), .ZN(n165) );
  OAI22_X1 U402 ( .A1(n372), .A2(n353), .B1(n357), .B2(n95), .ZN(n167) );
  OAI22_X1 U403 ( .A1(n372), .A2(n352), .B1(n357), .B2(n94), .ZN(n169) );
  OAI22_X1 U404 ( .A1(n371), .A2(n351), .B1(n360), .B2(n93), .ZN(n171) );
  OAI21_X1 U405 ( .B1(n149), .B2(EN0_int), .A(n303), .ZN(n245) );
  NAND2_X1 U406 ( .A1(IRAM_DATA[12]), .A2(EN0_int), .ZN(n303) );
  OAI21_X1 U407 ( .B1(n151), .B2(EN0_int), .A(n301), .ZN(n247) );
  NAND2_X1 U408 ( .A1(IRAM_DATA[10]), .A2(n356), .ZN(n301) );
  OAI21_X1 U409 ( .B1(n152), .B2(EN0_int), .A(n300), .ZN(n248) );
  NAND2_X1 U410 ( .A1(IRAM_DATA[9]), .A2(n356), .ZN(n300) );
  OAI21_X1 U411 ( .B1(n153), .B2(EN0_int), .A(n299), .ZN(n249) );
  NAND2_X1 U412 ( .A1(IRAM_DATA[8]), .A2(n356), .ZN(n299) );
  OAI21_X1 U413 ( .B1(n155), .B2(EN0_int), .A(n297), .ZN(n251) );
  NAND2_X1 U414 ( .A1(IRAM_DATA[6]), .A2(n356), .ZN(n297) );
  OAI21_X1 U415 ( .B1(n156), .B2(EN0_int), .A(n296), .ZN(n252) );
  NAND2_X1 U416 ( .A1(IRAM_DATA[5]), .A2(EN0_int), .ZN(n296) );
  OAI21_X1 U417 ( .B1(n158), .B2(EN0_int), .A(n294), .ZN(n254) );
  NAND2_X1 U418 ( .A1(IRAM_DATA[3]), .A2(EN0_int), .ZN(n294) );
  OAI21_X1 U419 ( .B1(n159), .B2(EN0_int), .A(n293), .ZN(n255) );
  NAND2_X1 U420 ( .A1(IRAM_DATA[2]), .A2(EN0_int), .ZN(n293) );
  OAI21_X1 U421 ( .B1(n130), .B2(n358), .A(n322), .ZN(n226) );
  NAND2_X1 U422 ( .A1(IRAM_DATA[31]), .A2(n356), .ZN(n322) );
  OAI21_X1 U423 ( .B1(n131), .B2(n360), .A(n321), .ZN(n227) );
  NAND2_X1 U424 ( .A1(IRAM_DATA[30]), .A2(n356), .ZN(n321) );
  OAI21_X1 U425 ( .B1(n132), .B2(n358), .A(n320), .ZN(n228) );
  NAND2_X1 U426 ( .A1(IRAM_DATA[29]), .A2(n356), .ZN(n320) );
  OAI21_X1 U427 ( .B1(n133), .B2(n358), .A(n319), .ZN(n229) );
  NAND2_X1 U428 ( .A1(IRAM_DATA[28]), .A2(n356), .ZN(n319) );
  OAI21_X1 U429 ( .B1(n134), .B2(n359), .A(n318), .ZN(n230) );
  NAND2_X1 U430 ( .A1(IRAM_DATA[27]), .A2(n356), .ZN(n318) );
  OAI21_X1 U431 ( .B1(n135), .B2(n358), .A(n317), .ZN(n231) );
  NAND2_X1 U432 ( .A1(IRAM_DATA[26]), .A2(EN0_int), .ZN(n317) );
  OAI21_X1 U433 ( .B1(n136), .B2(n357), .A(n316), .ZN(n232) );
  NAND2_X1 U434 ( .A1(IRAM_DATA[25]), .A2(n356), .ZN(n316) );
  OAI21_X1 U435 ( .B1(n137), .B2(n360), .A(n315), .ZN(n233) );
  NAND2_X1 U436 ( .A1(IRAM_DATA[24]), .A2(EN0_int), .ZN(n315) );
  OAI21_X1 U437 ( .B1(n138), .B2(n358), .A(n314), .ZN(n234) );
  NAND2_X1 U438 ( .A1(IRAM_DATA[23]), .A2(EN0_int), .ZN(n314) );
  OAI21_X1 U439 ( .B1(n139), .B2(n359), .A(n313), .ZN(n235) );
  NAND2_X1 U440 ( .A1(IRAM_DATA[22]), .A2(n356), .ZN(n313) );
  OAI21_X1 U441 ( .B1(n140), .B2(n357), .A(n312), .ZN(n236) );
  NAND2_X1 U442 ( .A1(IRAM_DATA[21]), .A2(n356), .ZN(n312) );
  OAI21_X1 U443 ( .B1(n141), .B2(n358), .A(n311), .ZN(n237) );
  NAND2_X1 U444 ( .A1(IRAM_DATA[20]), .A2(EN0_int), .ZN(n311) );
  OAI21_X1 U445 ( .B1(n142), .B2(EN0_int), .A(n310), .ZN(n238) );
  NAND2_X1 U446 ( .A1(IRAM_DATA[19]), .A2(n356), .ZN(n310) );
  OAI21_X1 U447 ( .B1(n143), .B2(n359), .A(n309), .ZN(n239) );
  NAND2_X1 U448 ( .A1(IRAM_DATA[18]), .A2(EN0_int), .ZN(n309) );
  OAI21_X1 U449 ( .B1(n144), .B2(n356), .A(n308), .ZN(n240) );
  NAND2_X1 U450 ( .A1(IRAM_DATA[17]), .A2(EN0_int), .ZN(n308) );
  OAI21_X1 U451 ( .B1(n145), .B2(n358), .A(n307), .ZN(n241) );
  NAND2_X1 U452 ( .A1(IRAM_DATA[16]), .A2(EN0_int), .ZN(n307) );
  OAI21_X1 U453 ( .B1(n146), .B2(n358), .A(n306), .ZN(n242) );
  NAND2_X1 U454 ( .A1(IRAM_DATA[15]), .A2(EN0_int), .ZN(n306) );
  OAI21_X1 U455 ( .B1(n147), .B2(n358), .A(n305), .ZN(n243) );
  NAND2_X1 U456 ( .A1(IRAM_DATA[14]), .A2(n356), .ZN(n305) );
  OAI21_X1 U457 ( .B1(n148), .B2(n358), .A(n304), .ZN(n244) );
  NAND2_X1 U458 ( .A1(IRAM_DATA[13]), .A2(n356), .ZN(n304) );
  OAI21_X1 U459 ( .B1(n150), .B2(n358), .A(n302), .ZN(n246) );
  NAND2_X1 U460 ( .A1(IRAM_DATA[11]), .A2(n356), .ZN(n302) );
  OAI21_X1 U461 ( .B1(n154), .B2(n358), .A(n298), .ZN(n250) );
  NAND2_X1 U462 ( .A1(IRAM_DATA[7]), .A2(n356), .ZN(n298) );
  OAI21_X1 U463 ( .B1(n157), .B2(n358), .A(n295), .ZN(n253) );
  NAND2_X1 U464 ( .A1(IRAM_DATA[4]), .A2(EN0_int), .ZN(n295) );
  OAI21_X1 U465 ( .B1(n160), .B2(n358), .A(n292), .ZN(n256) );
  NAND2_X1 U466 ( .A1(IRAM_DATA[1]), .A2(EN0_int), .ZN(n292) );
  OAI21_X1 U467 ( .B1(n161), .B2(n358), .A(n291), .ZN(n257) );
  NAND2_X1 U468 ( .A1(IRAM_DATA[0]), .A2(n356), .ZN(n291) );
  BUF_X1 U469 ( .A(EN0_int), .Z(n356) );
  INV_X1 U470 ( .A(pc_out_i[31]), .ZN(n355) );
  INV_X1 U471 ( .A(pc_out_i[30]), .ZN(n354) );
  INV_X1 U472 ( .A(pc_out_i[29]), .ZN(n353) );
  INV_X1 U473 ( .A(pc_out_i[28]), .ZN(n352) );
  INV_X1 U474 ( .A(pc_out_i[27]), .ZN(n351) );
  OAI22_X1 U475 ( .A1(n371), .A2(n350), .B1(n358), .B2(n92), .ZN(n173) );
  INV_X1 U476 ( .A(pc_out_i[25]), .ZN(n349) );
  INV_X1 U477 ( .A(pc_out_i[24]), .ZN(n348) );
  INV_X1 U478 ( .A(pc_out_i[23]), .ZN(n347) );
  INV_X1 U479 ( .A(pc_out_i[22]), .ZN(n346) );
  INV_X1 U480 ( .A(pc_out_i[21]), .ZN(n345) );
  INV_X1 U481 ( .A(pc_out_i[20]), .ZN(n344) );
  INV_X1 U482 ( .A(pc_out_i[19]), .ZN(n343) );
  INV_X1 U483 ( .A(pc_out_i[18]), .ZN(n342) );
  INV_X1 U484 ( .A(pc_out_i[17]), .ZN(n341) );
  INV_X1 U485 ( .A(pc_out_i[16]), .ZN(n340) );
  INV_X1 U486 ( .A(pc_out_i[26]), .ZN(n350) );
  INV_X1 U487 ( .A(pc_out_i[15]), .ZN(n339) );
  INV_X1 U488 ( .A(pc_out_i[14]), .ZN(n338) );
  INV_X1 U489 ( .A(pc_out_i[13]), .ZN(n337) );
  INV_X1 U490 ( .A(pc_out_i[12]), .ZN(n336) );
  INV_X1 U491 ( .A(pc_out_i[11]), .ZN(n335) );
  INV_X1 U492 ( .A(pc_out_i[10]), .ZN(n334) );
  INV_X1 U493 ( .A(pc_out_i[9]), .ZN(n333) );
  INV_X1 U494 ( .A(pc_out_i[8]), .ZN(n332) );
  INV_X1 U495 ( .A(pc_out_i[7]), .ZN(n331) );
  INV_X1 U496 ( .A(pc_out_i[6]), .ZN(n330) );
  INV_X1 U497 ( .A(pc_out_i[5]), .ZN(n329) );
  INV_X1 U498 ( .A(pc_out_i[4]), .ZN(n328) );
  INV_X1 U499 ( .A(pc_out_i[3]), .ZN(n327) );
  INV_X1 U500 ( .A(pc_out_i[2]), .ZN(n326) );
  INV_X1 U501 ( .A(pc_out_i[1]), .ZN(n325) );
  INV_X1 U502 ( .A(pc_out_i[0]), .ZN(n324) );
  BUF_X1 U503 ( .A(RST), .Z(n376) );
  INV_X1 U504 ( .A(n374), .ZN(n357) );
  CLKBUF_X1 U505 ( .A(RST), .Z(n377) );
  CLKBUF_X1 U506 ( .A(RST), .Z(n378) );
  CLKBUF_X1 U507 ( .A(RST), .Z(n379) );
  CLKBUF_X1 U508 ( .A(RST), .Z(n380) );
  CLKBUF_X1 U509 ( .A(RST), .Z(n381) );
  CLKBUF_X1 U510 ( .A(RST), .Z(n382) );
endmodule

