library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.all;

entity dlx is
  port(
    clock
  );
end entity; -- end dlx

architecture structural of dlx is



begin



end architecture; -- end structural
